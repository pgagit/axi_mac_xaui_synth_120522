`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
B9c5dA/oU443B3GLQbhtxg2NW+1aJRSo0dL124shpSSz2qyWdtIYllJyJOBbxxzLhVQHru94Xahf
rKUFgUsXeA==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
e3JD3aoQIBAsK3re9WaB05Az1N1xrJwCX1kJuh0zu16RBTRn8mmoWnAibrnifCxWiUm0c18VQYKX
4hUs6BECXYR+IWEy3Klt2twozDnHdk5E27r8V6unC5VU7J6f4cLEH0sw3iH48lML/WXEDlq7Udai
IKh2MdxpLr4rxRczOGc=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bnMitQjc83FQdVMBo1NkM/kItPc2uiRW/FIjGy6R2xiGAC3qeis62RHlRSIK/i425Mt0bfN9GSyp
st5KHYxuW+Ef1uNaaZy7s4GgrPUuRsXDP7bHbsBcZyDwoDtTgYovhrERncAR6EfG85MXdx1ORScJ
KXNzLa5HGVCJaiiT8gfVQSqaq7ztNWy0f6PCYrWFtVBwwpF8AD/YMbK4VeEKvMCIoXkvn6SbsUbR
j6HDCbyeIkqhbq7Mf1sKbn7bIWYlMUUscPL8nGzWQqTMbi+Wfxvj/caDJefLdJVEvcKXqYL2u1qa
RLp0QU4mrcN1Hs3m32G0Ce6z0WVN7XylSn+Bsw==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rS4XWuq5DhqyI4gzqNtzW+QMYXOAwcgxeustSnVfgkpJgD1agBQS2BpJJ1AHLFE+/RFpBY2pSFio
siO/2rPEyG71eUDu5BTf9zheuznUJ8iE+KfFb2y8VSpEbasv0RG85BazArMJUJ7eC22j70qo7fSv
s5oRzwo0hueXwLkWmXe0oipfI9mWhSTZMcUZNJx62481jpVVfNKPS6W8lffAXm+3i15HFuaCDYW4
+1VT2KySKtN+VIrz0l6NG3lrJfB+tlFPkvJGRBvlhTzLLd08ET8uXGCvoeSuG6O5OGcC2Kgg3Puh
k4FRMF8waauEU93cfv5eyvuix1MfMngFTnCWbw==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
PrHDJuzh5zI6jvZ56j7/SecSi83niBHxd6xpJ92/XQQ+AFk8FN3tYTrRElFqphcnEPEixk2gwB32
/WofxDs5tydePqjJHGYTytle53Xb6YWDJ7Y/q2f5/aP00uDIYJobCIMo6FIKVWfV5Tw417eySloj
6r36SZ/EXEqt4UFBS2dmC8mNYtejPGP9uXOfhEimJn2VaIY+wKT6XEveibEFPhm62ssxVpx/Kruo
ttQtFsql09STXsS63XdCGsmBl3jyiZZPrGEWcHsyvEbbtjTMBWwjeRxry2gg/ErvyRsOEV5xOuoX
e9YR88ycLLizTWl22pGs4TASwvXtDcg46nDwYw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
YBwqnIpw2YaKpW9xXGm8s3qz4QphZdTkpadrj1GFroPPFT9InvjFPm/KQZfeSOtTPqiG51Ped7D7
WP8XqJG42ECjG7z9pyaOWMkKFFIM24SWtBeWXLYDpIzQkyfo5Y9fI2++08CRckiW9PMEdA5rZky9
A8HnPLcarqo2k4eKfIY=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
RdpyS1Ye/C0E5kdTEb3Af9+Kk3puQlgywID5PYihfG5+uYwURKv0Gde+XodAdx27tUERCb8B0Ftb
yDrZsLWkpMXKT1BFtEyYpcymjBEd5hFJUWJbM/QY3CD68+7szdv/3XrueC+DTrnaMN5eTIdPmYo6
xEC3q9ssAnQjS62C95Dmr861KPhHftB/PPCsUWpJAHn50A5PPvIybibh4roE7BZo6rtiDJwFz8NV
LHMFBGDxH7/q4cZG/a5S7HURdAsVgjQZmSfHijK/NO6DXhsmn0aqbzOUurrOQJ5QxDpEeaetqxiM
InpA4aCsmCWaqwpX/AD9JKyCqprrCCD409K14A==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 211040)
`protect data_block
n72CGV7SUiciUNjxxQT1WzyjjCA2wJtqnVlhstFDayrmuDmS3tE4Hg+flGCJ9qUSOUkL6dLvtzCa
JIQLsyC16X0SRSXjf1J2wu9kvyV2H6cN8xb2WMbxOkvGwY1OkXbKSStZMIJIwaTP31ApE7r+Oyry
gHwYg0bMAUlyMJs2SoFQJzdVozYbQzQlfEsr05eYHcsOmF3Bqo370nWqWVb7pnaA3UQaGuiuPVWd
3BZXAE4NLQ9QdD3TF5b5NseaNP9MOGO5btx866FupSGNlZ+h4+VfCGFH+hithJiF9jgMw+Vs/o5I
dyr+oBZ2+p5WTl/1ovekgFC/fDrIQOlBl7/migphxjs5EmMll7fU10+3BC6+BD2phj7CQLG88vYb
yi8GtQEjvroBjVDgEY1zWoeE1dEyoCaaLW41Tqu0CYHeRfGpjHi1X//ZKaFbRcNKe9FpiN281EPc
mN50hs1vA/u6sRXNL78cwNhMRZayL7MZQBAlHJCeMcVl5Q65UFpTAitgE67LM2wUBrAuvrmw4MJF
9YA327LEplxhNqaEmKYbLsDyAqxVYqqpd5+7z0hfYc4GZFKpuesDvIqzWZll9UYisF5G4DRTB63U
wlCKnELJn0uD1yb1oQJ9YxzAGdQgcmbj7Ms+cn2guzIc6YFEjZkqPX0RlDBIpGl/tz8eOra8obvV
AwyYHRqIg5ANBw1wmjKGpdEkA0wtPkqkju9gHHyN2wlnS24MFDAofphtDJEAPyJMy2odf8zizaN4
oNAsTLVt9IGrHDLTJ3CVpiXZa3hHxla6EyOddjP2hUNHOz4t6ckFusHXfC9Jk/G8hTto1LvA2Jq8
hU+ti5HAZdSJ+eOkSmSnIrmKFithJusLLQ6gaL7QNNq0zjNl87QA7VDaC7sikvfT3ICzQrr0lqUH
HfJOJoz7n2+g/SGf07kN9axKPPGi3nfavJqe92iZlqb3uVKPNgyPJbbsKKPJpIi5C5p8cGAXeco0
Xw3uQvJNAU4bSimJGHnGxaUGPoYr3A1aThTxkbQi12GgwmhLJaZCxBEJ387aOPIAF0uCEtJ+NlZ4
gHkKOZXbYpDOczrM4XO5dn5Xua744SHDH+hkF1GAPX+KQfXy5WTLquxSwy9Q3PI6qcFrfaj3Qpvt
C4SmqkZWdLRlvRCW2q4qrF4ld2GCmec2C6iz6bTzo67+9wLZJ0w9dvETIm4mdcd02w757ChjKcaH
65PJLlExcog8h2b/qwBINZKulrEFUf0S1NT2L39eKjQoVtICzUE3JUzecc8/dupTI6DZcBoICJxp
Myjh25Lqs0oqo9GfQZfviNE9yISJWkGAq1/fDifKN9WtBn4sjXIqrA1IxK7dAMFtIHT6oyORoBwU
JjjIOIy7dhC50cbHzANuwhjpkpecsG1yqbKxZ/Wtr0/mynEp8oVDv92+scjfANvNeb4vcHcCDKDn
eEOXhhoV5+5UPz0gF2oM2CQUGqRvhs9av8MGna+pWC8BHUueG5kdIZiSPpkiI4Pc7edjMYcQ6WlU
2T2m2bn2cFAcmztfzcaQ2OcibBgDwMoQEHVjRstDlU/0cMIRLUGyPLOi8lhjXoafP+LcmETyuTXh
my7bLJPCaN/iV04tgsb/54H4vGmVKS/UGCaZzEoeWgKpAmDWB/0brR1xypEUoR20dyXKe8FypBgb
6XyEGG9hudNATqDSHM0e6CJHXAr68F5LSygbxr+60L8bUQQW+ug1J6Fyii8uKWpcH6NLiiTv9yJ+
YbE+hCk7Nv9v29xJU/elmum9IiAysAh13d81VfijMpiWc/23UIYlqxtO2xosR2lqPYglq3nPv5dR
lzEqgV2Lplsis08oMfW2LJuYH/lnA69mBikDDTTFfOXFDhQVoAYxJp4gurVI02w3qnxbcLcoylof
GFHUVgWzNcB7swRwNEZV6CeKuq1+sX7jXKP8aJENXyoz3vnCIiKN8a15JcrSbIyf9/oOq5hcwvB6
DlwHcVyoBd4ty5PAUzN85n6VZT2wOfC+9XPAWpq+SQoF4i230g8dzGvhMwDj1BHBn26hokvop4q3
vSA58EB3mJgIsID4/YAQa0HYXAI78Uw5ACDK+GPfYgjgq6CHb/uitufGPCW8LNdogpDBjj6wlxi9
iREuO85Q7gXGU9Cxojf1jq7J2KnrH7Q4w6NHxxQvcwcw0Fopfn0wNKAwiNu5UKryAMSOjJwivDNV
6ZK7hL/cT2UxgJ3x/6gk+swCmAQnVez2+HuyJEiMNxU2/eYgBWXtA3DOHbkjGiLpsUHXN2EYb3DB
gLbMRX9vP5wj/d4M73CuRUExYG6wWakLtoGWg90Eg9n0WcK76LUjH8mtT6zGRS2b+SQvpv/1qXag
krg4D9yIAB0Lp8abf/nOFPtWSgHKiFkMhrcvxNtB0FbnBizHVrXvxrZ8G8gthL6z7lT49bzlcoSz
b1K6KrzzCsDm+ODdqK4r0TvKxaL1q9XScD0IBmTKnI2mPX8Xkh2GXJ9aKaZsK4B+QFR7VaVzodN0
LTkDu/b4oVn+8yZbejAfO6eGnWtZPCgoy/iNhsWpz7agqfeZv3FMEqdentXkI6ueAe3tXWvRkxNy
4OQSTYnShBkCr6/PtgawNoVT9KMthJ5gNq33DcVlQwMFJtqhLP2m7BAkyp7tn/AQ0MEzQbKr4qih
pn9A7/xjphzUZRlkN1n0nejYQUDhJbjncrVVL6G7Q1r6xGuIVfKHBjou6EC8m152z6FC5lAQ9Vna
5NrtXLSOqTizAJeajwvjcQYTUi3UT0Yj5lqrWhDLj928N6Qz92ggk5d4RoARSlbFRN5f2z+ENGus
HyrMvClDQmHef1+qtyIJPiB7q2blPzHmEjeE7XnaqYTkqtLpwIVH2O+Ne0feRnSqewTdc/hrsYLQ
m7grpzE1yx3pHMXnUE49i+eKmqEppyIosph+bFGgmPEV03V0fgiX5uRUAJiOHNytrAysa7f2Blk9
o+31BzXcjhXYG9tk3SQJYNojFvH2r3N4L7apNH0IREka94HQ/19oBhkHLZ8XXEoFvFzyFektX5Q4
HOZBvYm41E5nlB0I5tzSzupWMX6saolczaGKeqZ1095YCej81veqm6e56LHBvygNsLjADTbiDmKS
v6XmlhGdUq+eWv4kqLa2NDVtAUqjXUNirQUWTUxnz0eWpdqwGES7Ymtytb/0SoN87SjepkVfalMM
vSMhhAaEGdPJ1Ov14/n/B3aOLyvq91cydMDVOebY2JCsU4SBdA/5QWsl0QEJrezvOLD6XI34RpZ1
6ZDgl722m9+IahVUzoqGhzcDHZQj68nHpAJL0bMvkm+GpRtESRUCVp4QyPhdPqCQ5UkDjROYP8lA
7+s3NY4tJRALAaT6pmbF1vb1QWCg3lwGngt/kZoXTrwGONMjsusW+BseBC4MoKtQeRgBSxeRyR4X
pDHPvkb1D2kbM+5g3uszS1izHzd2RyIIe/hzx/9KT+5u1ePYLipyUEmKf2/RdDWroXBrU6SDyI0G
Lb3u65SNyuWEozXqlrB4OideepE+xdS1sz7bx8eONHZsmACc8Wvh9stvUPc2G1ufXesIDBLkNQoZ
dS6ymzPB6+1Ye/BQFj0aDEHnCoEgvwEe2nvwQXKlPTonYfEeojJ/seuQnPbokvELvDrFpK4T4cWe
353ntuqMa/Z76Wm+fGdzsBXbZujMqTCqB2fBDX554Ac9UUTEy3sPwWK0Vz8yUYDtJy33jUgtmLLo
vLjLvhFyXtuyFiR2YNHPQfrONzVtiqBTqXylIRwqR7zy4kBDBJHPbZvEiIVcxIDEjZKI4e5viVXp
cQHvrM+pEd+gtw3JIV6srgsPhEsICidyPmS6BWSw83jp86SJFjWwEZF/TfbaDQM6Kp5VE4dD1fxC
PS9k3/6S0isbPdo/oUiUJjznXcZNEd8w5SZ8Oi8W4ta9LgM03Zp9DeffLRIE0oSog8d45zkujpAQ
Y5dK8FXbrqb8yc1PbQQPr99Nc8+kB0u1LkvUA+71J6BcfJeX5OrC4GqWqeyn2pVBH6Q7EGa3arbg
TGS+pcZ4LSf/q5tAF8ZqZYJcipoV/cLGhupDRxBYW2mhRVQTErUVGNtsuGIRECiGDWoLG9Il7S/V
WSukmpObASRInapjhsJJj9o9V5BY0qfhR5DsH9T6hPUsG4o9JFMPSfhvuatf9HqEBd0haOvisOKJ
VTNa/dzQpj4/U90gGp7Hpenc2VbV44uhp9Y4w9wycSFBs75Y7lfR5qmvsZx4POsAm1SWFptwRxUo
d3Yto6/tpWBcc4bkWgRLX1ry0GwyMIISBbmYOQsIkulMtBMZXtI5eWkzLMXzf/DpE3XJBeoKbpCF
l83GojOJ9caiwyJw+Rro9Lngi4rPatat4qTq8O6SQHNcT2+/wERvNOK6FBKw2LSGO+Zuezn9CmNd
KsEmuL2VvLdTTfQG7e69VOa4yV7TYjW9jI9u/IWRNef+4cqiGxCehs91DLKpLRQCCjoiF3EfSLw5
8id52y2XA4eKXJeRG9G7nxymMqgL4fq+r79JeWYJNiRxrzb/cmjXN5dYnVxgTjnTfKj5atDwTn5V
TT0ZkMM4pxe7w4QoSy65928K5vpsNarn4wvZO1isZpaP2rReB5A0gshHPk+8shn8kZ1dW3o3qty3
oNcL6/2NXOhO9w8sAAhMMHJ5LFJ7QWqCoYuK6sqsKbxf5iyk02As7EQoI0ubzeFSKuYuSrhy/Qg8
mbNfAZcC2JuUh0W1GlS0KG70sayTZ88v3oIbTN8LXeYUdKWwBNcfPWLpVJpF17vtbu0JWwzYLWMo
aOIperc1K0NJPtZLdEK9tQqECUAPq1ybsEKQcrYjZwFN5h6q9sLooLVEeaUa5DIKbiO6PwJnG2lZ
l/QOth4Im0ducdvTBdGefDN17FfZCfp4Z3/c5nxevygAHebFia5hFGWalHk8XYp+e/W5iponnmx/
/i5lijlNW0Dz7+rXjenRMsgqr7WOkudN5/CvFFZOlNlhecZbidRxfemGetlsaK1gVYQlB1n26buE
BAg8loErTl49XxLaQk6XfJid6B89FSSYXCAEhoqqPP3uLb5c5dbU3dLUbh/2gxek8tpFE4iW/9ua
lvw4Xp6CxkoI2p+Q/XasKZeFKYpes7lE7+3ScPgy8DROmkwFd8QHacpAEtTVPpFShcBFgDJ7gDCc
gxq1Wd0zSo/sO5Ouh4INYd1j1DAyli6gOZFXcScQMgDJF+m1xYarm2mXq86VM2DsuPjjsdYnpF7w
uBaxidO0Ct6TTHhysPBHJvL6W2ZDy9tJn76W3yu43+IWxcq+fUrhJS0vuEzQDocHpug6mgpt7V/J
Scb4CRwBBcw/dyvx1chPMrIeK8+MhCDU+wkLJgkDGMkoIcV+SQ0NxjEgOsNYXCsDwkHZeAxTN9Re
nQl08VJdx8LrWP2OVwSbwyhaUV9uY+eUcGgPpURqxFuCYECoqwbV5gaFuIH5Va8T5gkMPS0S1G9U
fodCSogryea0Nvdm8C9MIKo3GILqCDPOakNStcwONf77IXMi4GkO9dyEkc7D7LPOueowq3gk4emJ
2jJXFdiZGi7ZRMrzrR9BlnTSHom/S86UIISAodUxQrqCfDY9WLXZt7FbxZmHNJM8g0Dh3vBXKsSw
58MiwHMssjyPvLQ/zrN5x4b642wstToG7DE5MkpQYKfJ6JWr7WLc2vSIie7AKmc8Q+ej2ZPNWlf7
ngE6XZxEjpHQseGg0mq9lHD6IG+tf9wV1yFmJKLelfvM3y9K16ET2cHctrmW9tZ/PgpvWY14ln7C
InL4J/KWUc7WNYCfdGaZVrnVmponv2X+p2tM/BhriVBtabQX5PFfmEwbETYOFoMD4Sr5x+4bY1fV
k2hRlElYvL88u84q2X8QS7RQvGYKl4+0lgT5Sd5SvQvOAeglQZBL4+s6ZlDDOFf8Wn9a44rNCNOz
fVa9K6QL9ePgEhIi/Mm4ZRmpZg+eQry2j8Nz9RXbWpmbqfZgfnnNPhDHB16sGTVlk+TCIjwwArgf
2gUFmP0VRmy7vJShz64jpMgzQSg8BN/a/P2HHBLwvHrBRaLBBcgef56qG6EmTxWMRKna+9t27ClW
g3IiiBZK0C6hrS9KGvImAuylsFsFyVzC8V+50slRY3Te/sJMkKbE1j7ntWAQwhRP7MOj7U4epL4J
oaD5iWyIyF4eZbMC6m5sR6vxGgVMLdQxOwtUh606lEgy0vprFQ8D2Y4bAeWaTQPDux2U4GYlBhBD
TZyTIMEpcnaZWdEPm0LsJpr3GfDtjeCHE5wVpiH3xr/4TsWS0w9XJ8Yw1hcfnrbfXEHqLrPXtFFT
byj8eizQLsG4hYVY8p+KsMvlcnOZnINK4IkzyI1gpb4FO4abw+0W3KFSI6R8ZDwGJjiauNY93Nh8
jhvPkZdM2U1d5SCoLCJNFKkcf8zuBHtssGZgCc42tSNnrMBXAzuTRy/bBRs9FYeffdWgk/yo/4EX
kws1ll/rCBmLfxga/iDv8rD7B8HArUqLl3ZesJ7xSri6t2OAPNYwfrX17ynbmZmEfHP3rDS/F0xC
AiMdIl1emp8QcCuZVpOplMHOBl+R34QloD33UxlcwcYP9LUA+68rgUBb9Pq4rCNePg+rh1yP2COW
/0xLKbWox/JAJD1bghN8Vg8VwtOq5GpPkb5ltqA9eM+clceVI7AezyAFv/kQBJPzbi2Lxl7jbh5F
NkIEWFO5+iQ4dTAqE+zze1rWAVJFN7SvPjiWrgQ2N16e/pGa9pjc+40z5/UH0/z+mJM+HCrppSdT
rSrDrJwo/mUMzc8mbUh+EdXGzS8pmKYZvGUxBwPtr0fRQrta+kLyeF2va8gWUh6FAwPMjZQI5NXq
HMkWXPJSD6x3gAZ7hSjNMXbG2XZQQTUD3dLM9m21ytyv79VdAzUwzgHCqI9nBdDVftDkGli+sQDi
d6Wh5GIme2XKZG41Mdg6wjMFYWQ/DingHadlY2TWdDT5TK1RB/2kVBfRmO4w/4VzaVCdPB6FjznT
l3qgsPBPLDm8JvodMmG7biUZV5aD3hB8shNpF2VjFITllYV49UImZLkOAtaqkwyODmellt9tQlB/
QfwCubD4zNE8T2NIKfU4f9KI8zFJR5m1FhCghM12MG+kkHzR6vgLi/Eg5vQ9JQ7Pe/I+kAUTgd/9
H87sVF3JF1o55X89m/ux/IlKzJMhLOCkNiC1U5q43N2pTScCMw+AIAkh5MGoUXmUlk9+AX1nWNht
1B2BS+pzjb8D2IU7BeaToaDdKWSmAtnO6RfQnyZBX7Odlz/MLiSOmncSxJA12/N1KT3rwNyHLC9Y
PfRyhn4PX2BxPiajWiW869SqSNyKLC3oMJ5GeaqePAJtDppO3Y8UvIqyGYBmMJhGJDRhpo+sfxVx
gBXPyOO23Gem5ckmOyqyod0hF5ir/pM1Z6zpSpDANyAwRWkjDYIDAMizR3EoX8chx7XdSSBD7O2O
0dmAOmMxXWy+/y1g05e39T7QFIojtAFVKhBMfEwwa9RLX8oty/VuJXXH5YevzZiwnQSGVpeUj8i0
2SrZ/hEK6IZtYh+0GuBteQyOg9koymZdzc+/Cv1K6wX0O2NOvhP/OgzU5AJXC/dTOQ+JrSwCgyeV
hrbqbIMXTkSZxiubBXmXG9iJ02suDdvYdg0IBxDJXL3nJEgvDUMCOgQV1MtC8u2RYWvsqvdCG2uT
88eZt3yGsLyGpVTnyjELOiNJsVRvKjzcTMR0clWcpMmzWiA3hAtTEca4rxW50vI2e/vnqjh/ghW7
Hv1k8II13RvArI1GU7JJAVFqdmgi7r2SROlApAo9Ciz382udX539A3n1Y5mvomQmSkw2mZj4UoHb
vgcwA6cvtW3z6660R7pT4gIi5uhG2XpKTtXZZ1K/GvC2L7qp7a+J3iIcQIurVOrkMWnE2tKNhkpq
URbfjur/4mcO/H65KxwmhyCAl4VHy0tOQ9DqREtgn9xAIaiw9z4qjFm6yGDCRjuKUk0mamIZYScx
xHehlE4Tin9a5QOq435KCTNSgdfWLu3Wqc5zLTwwY1NOke7qTwZUDObiECSsLeUwMLMHU5Pqt6em
q5CkG5N6knx0CCuuQoISahLHt+RAfqzJtbzrhczdOeUqroywjwz5apV4iL1ks1w+URQ5czMBkz7/
pnLCbNStg4PK+qHp0cSAlNarE/pMzYAFxqwKEosP5RnjADl8IsrywgM3ZIS4BB5jMXoNZKLLnq7s
HO2NcmB/WRI7wkis2iR196z31jNNqJUd88cgLx8L1tEbt/x+8dMhTxp6TKsHEthUDQ3ESBaQR3ds
flnqncmsgAcIQBqNuzIR7uxjtjUVc13fSYMWLZ+IInQGvTVBDJXH1cSzkXMmM04J0J0euoI1LEhh
g+CUA9dModsN/SHfXfRSFs2kZgxwBuNIXc1O3tkdwUybwnrV5k8YoP4JdkelAwGoSHLvDil765EP
OcxWTxBW7ewm47Eln7hgOLEePtP11d4NGfshkQZIYQGNDZebH5MaLwZorNlHhAMu2UQDuvKJCKVY
8tpAaXUNpO5zldMTiwXh/vW0ZtI77nuLicbi8irW/sNySRQ39fDKuqUG4MxJcydQhy00C0raW/2H
F5zgyrw2p3Hc97H602ZXkOsGNBLqBwHn2O6taVhTW2snbIMwBqyIU5Dax9PXO1gra7CV4OSJHmtO
bbVNJaI+ZX9wQ7xGSi29x4LTv0Ot/sgUp6vROTDQVotjaS8OFjb2+fLILctbqHUGoeYtmEb1Vfes
yMHth86mS6WtADua+m3o+3K7CTTe1vDFJ6Gs87/XGd70hKaFndtQ8Ra9WqSAi3cKPl4g+zMIiM+2
3yaWcI483qVdzG8yrLISyofKLDzYGZxQagUxlmsqIEuMVz8x1LTMhOgCR/OYdbmIt8e6rEPYabJO
HrN0KeZXe3dpIHoeA1V2lKgfe0uEIuZ+W2H5AFAN1dim0WEUCpsCVXehT1dwUOx2YPazp3tvnDQ8
xRCIgbmhOLq+ZOTpRSdz3FtlDO5v5h8ueli7BJR/qOkKXKndRdv2lupXL1sUcsB8B7FJXL4eO/2Q
Km8EASXRGi+UeFbN2t2LYMReR94uVKB0V7Nc4josbzaA+nxdlwkr/QS9nrXGO6dOmyCOLax8VDXg
TTTeP+lbebcHkYQfmsAAQEYC5FKYNcEtCIM/psqyVISIAxSbLYLeRJWrrz9zppXRCO04tm3FTbUf
Ep/vOIlgTleyV3jMWcUuWLzedFmyK83AMASS0aq4j69PV6RA6A3v85/wct67lcxcR3td+lZUdFHv
sL2zKqurcCLSzEZNFTinLrcJtz44b9/uPw3CFDkCUhUMiusc7LtvjQnEO0a3XapHwLGBw3PSYBh7
87ySE29QHzlarB7YM1oLcQJV4w0WRODBEvU7l9nAPFIaIMrB5dsUvwXmql/tWN+g4rQw32nrPK80
goi+jlILlnYobtzdcBlLKMmcxxK5Movvu5n0cqaZVYN8QiYBkto7DfgkRs5B/RY/9QdeMcsXiJDQ
E2QdVaPX20jklVuRWlB8Iq96yO9TkvH6rVy0POlEMnphVlcZARAAAzXshv7+0g6v4DYjo1HQwUHS
V3EwLrFVlPi2cKvsVOk2rJdpnwjHVQVENWfUNoDLAsapJd114KA82seIMYCtrEDbtip7vFs1sWCP
PjPuJfHzjhJlUkR0yB1/nPAxufhVTjjcp2hU5WrLFHAnkHEC5/QncnKjJH31mqqwETS1IIlTQmG7
LMPJ1YVz5B34tQrd5wP+A5aUBbwbWhwgzst3d2StiAuKKMOg54eRUzNGs99J97V6QrisvNX6ZfaP
empNvfFXbHcUMEQBjUcrjTipElu3y1ZkxnJcMAYJjPPV27MO9kWy2K9KpxgUms3BFltaogCV8aFU
iAJ/q1NDXJ5Xpk6bS7qqfjacD41A60fBy/CMiacrhrh0OOVEAe79Z0G/ovT1lr5jkpKfhLVIyCYU
mVTVumxZULxXKBnaah53JpoIcu37rl90b5Gdgdg4C7WLsFDIZ7gHMtPJuzxAK4czNzxpBIN0H2bg
VMr3Pw0BJ2qPt2dHugdEcfw5xKhAe4PjF0RwgG5+QSw+fmmQfYKx5r+vvxmWF1lxmoZw8ksLVREi
JNjXZLugv5zkSTunudu9ZtRZfyugBigp1IPQhtwGMB4kTxDMpcIMp/n9QJ2FUz6c7R3E8OETk6Au
EVUnuax3nHo35VJfeL6wxcPLagkzXTsPbagcqtqBfmVDnA+AQ9gv+HMprGpWJw5m9jhNzUoOsF/1
KkOZ9h9Be29Ww7I6y6CCCn86Uu59CGsM+QqBYTP2D5Du4Q2LRW3nNYovmEqTvjiZ0jL7dIwD87PT
s5Z/b3zgQ69QOLpLADAiRdbmVELajJTjaQZ9z6sNR6cKhUuX2HzRmKnnye0rgKMFh3Ks2Uu0H7mc
CRSLrKx7zAIeM/R4FKwm5NGGRz5gyINhXOrONOdHBxG7CLMieC9wDeopfJiCnohVGuVJkbJa6eLJ
YPxzQs5laBR0jBQbarJBodAn5qg9q29i+hsEzPX+AWa8Fcdl7OSIZXrMcHun5vypCwwgDfeQ5IAN
TfvJYT83/GkcLdmC4Je5JRNu6yab2zYECNhIBujlGeCJ5AHKmVK1hhjDmMZAGLwIKaTN6x1ZOMNH
gdDkp7SWEMDZaFcO3BWFgxiGLzWK0p78qAhVqqhPC1HNsVyZliQqpy5JmvLf1AdoY9VhZLO0FTzM
kQJGScRSlSnQ7H0iUOR7ZAiGiYBLtDl1JgRIW4Z/mkpkysx5gv+9bDLzLQIeRL9xccr1sEfo73Eo
BaODT0rCjLUbzXFKdI6NsKCJUJKDHTZF5DCVw3cIY32rmXzy9i2DSvS6RZMkdQpO1Ao8IzYfxD73
nQFwXwa0jX0ZHbk7pjb3aF0/c+s7cNxl0u640wk4ZNiaHeL45yloMANV0zFL5N2MwJgY7/wKWwvL
Xg5ZBUPRMiwFBbZ+WhQCvaeX6OkFe8qcn5TQu2t+cPRnU+7E8ceOJPJbNYSbNA/M7hZWBekOQTVw
6Lx/O/2h+OS4CqMlu6ewcdu416/tzhK3tEmF1ZUt5c8rAtRUJei5IJ8GJ63/Fx3HdsS8UHvQDR71
Al5tQwB1Bu3lv9XG4Mibkm7bZT5/Pq+PIctEdE01A7BnUsIwUYNxRkhopvgRs0uVVoM2WDTNKw+v
Lq6Qob4WwZXY4MwnUBUOl9TU/JitWx1WRENkioKowdYB/gm9ZV2oHrBN7UqRXLw+obRmVqJXyfk3
/Kf14wDPPIHQZ9ao+lOR+vcSKpcu6kE9hGvRUoK+ZjWtEyEZ7pfGyf1Ys8d34cNCeB0fYor2eeC/
+23HWKQnhLxoqMDSwZrq7Cl+BUjg9/S/1JXs/8RKICNBihQ3HJVQjMlkH3kCaoGhIwFbnGCU9im5
KkKgtMt1koVi4SjEeSydKJL3VLSInr7wy05kEg9uuxu5IqZOKrye79Y7YHY/NiKlhbBjWhU0OYkQ
BdXKFX3A3gNxHeBISzlkRHDqZNVH2Eof7yf+aRwfqZP2StNdG8LOX32mYLGG4j7XjnCwdBV5wi06
zj/CT+uQnWdMZ+Jf0FWskAnsxb6A34HCTaWWdXiZ70K1SDHSKQb0V1oqLHVaPyXODiSDpjHcVs0u
O/UVQVQHmQuOLvbQZzZDN7V7OAZ3WTMvWFo+ET/7aEjr5n3Q8MRmD67o0VNW7+7ZAVW8D5liQ70M
tF3p3KlSee/Coysw2i/srV3JDBDZnmNLBh0yPT0iitcAZK2U3UJ9k8kiB2dwTa1y2Ub0XKPVnK0X
sSWhIs0xVgBU4BnHO2hfH5Wzip/b4haQmn2z9aZEPNR3lS/uFIf+8/1VOKpP2ymBU9ZdbFJC3psB
GS3qxlkqN3yTmBJiwWyIXldpUo3cNBwNbmj/zWFELnHT0D+YI9kV1yl/mUfJ+WLuMMcyrQuOHHX2
XpvyQ8qB7RW6yx2pdyvC9spnkluFPUMr7yIWn98dgW6f8l0RNtKmSCzNp6/vFcPUN574BXBzTrKE
Gdk25eS80Ffsmg/OC+mmpD9H0k3jp11TM5zJsG/2kkT6JS2Zcza1oaEiCeA9OGFVjP/WXvAnRWf9
3jBZz6PdpqKDXXuklDGfDseharf/ad+t3FL9ZLk66BhFlsU4ljnrvFqvKEHBfrYa9ykio7Bzpeai
tQugkH3IFvlBVfjR1tfi/cIW/VLRtGzprh9htJAvaMk1Fj9mbXOFpK8vUBSmyyaoco0niRBRbn+4
b5RxrYu5da7nQUdF1EfLVOvUoUKuiPyucV46kESEmgfnV7irz9etAwhX8khcQ8M5hrODS98h1VdJ
p9C0QwYF3balOy7l7842hTA+Q0cFh6q5S4MeDWi5JQ7fsZAZKcw8YVKyVJXnsOLsCD+sT11vcN6T
EybEZDSdpByLEd4D4Gc+lIDNNIzaakm9UJ9+Ofx9yZvb5llUri8zWf8SdACP6M5qs5bfAk45iiAP
Z8UnsHq7xNiNa1zbaX9vdQKaF43kQFuocMabiSxLim7XbkTp4HOi+vuzVkOkkUW0LyY0vKyeoL5V
1l0FKJJlKJCK4Ntj3Qs5e8IiuFPr2GG1KpUZgHMhJqWF7oqgpZaXrK1CFpd0vi94t0Rf6TGeLwQN
bzU4IAByxWfI9ZZAdVTnDOeiEFDJYr2ABms/Xn+zHoqiiTcsAx9tor+r/424FDMDIbbezyYXFyFa
uJvHEAP+UKM37IPhwqyDgz2qk5v0mbs/6K6Dv9+btEWlUJV54AixBCV2ykSW/7IV1ArQUesQr+Lx
eR5Wpwvvg0THttR4KIfTDJAju9FPkadRj9xtN/pnjp/B0QfMO3TGmIJFihhLXOQ9awd1JGwYGSJp
oTAg1GNnwcn3kq4hROc+EZq+dvKEArXCOe1mEW/Q4Wqz+4jgQ8paB/5ZmdwVrX9I0wX4h65e8leJ
ciWpcWsWwqpl8Pyi0AuqeGq9oSuxWhxImlxRKqj7P6QpLfCzulWKx8ReKCHjLtx/8P8iTqC48ggu
BbfT4QVi0tgv6IW0mO2qG33T1B+aPgZ7i6i8cG+mNJF1Z8AfGIbAdtsQNgim87f4iV+lyLI1XUyH
/0qzOb5XCPob2bc8IGo9rneKL0kdGybVXHcziEzMxgjf3FMHGO67eIMTe1Tkj3xthrcGNx+ADgib
3r13j8lh1zDs5OrXRbgs9PXtLYa9f18AhmGnMw8rvYJG4Ja1Fj2Mm6g7CgX7YLd5Y90D9BzM9wtC
jts8wJ+0CeTAGDsgbP9Mf+xqKXy4LVXm+srE6xKEW0KkW9Y1OPRw1jr8i/fXCXjEUFFn1DlxSfeO
YVs6NkUN4hR1Wx3d6DYnavrxvnfrvdKNcsvmDu1hvp4YsE/4F1NFfnv4K5+Nvfo8Ltg6ErC/aCQZ
p4dbZGtRm/2qXHQB55+E5eZaBvxV5QlYHX/esXJpEcyc4X++1i2gUIGtbZTaazFuZw2u/tyH61V6
uszqMuQSZHqmFWuQnrb+0CkwCNXb/5hgRZ8pKKEBlqdO4VIZKEbalBumTYe63v5r/MRDvVWC8hg8
Ki3m/0AGrhK6h18gnmwz1cGctJPBxONsG9FGZYqUZ21acWOu7MbfNkn/X1oeQrypqrb5AmYJkmwy
qLcXMwxfsweNj2g/nktXLPnE614Bar/23zC5eVGdGOyTVLbEWHW4ErDD/QPcY8ZzLcp9O0RZQpTR
HjtvF4o4dxg22Bz5xTAaoKNDqVjIQ5VpQQR18h/hG9R0Ff/57aUt8TvrVnSSJuhxH/ZVvqv/0t1k
uERbQXwnydLzuRBqGMXVi4ziVP1B9gpG9kWkOz6YJ+WLmjbtV/vUBxmkbva4KLAWwJ7OjUNeEHjW
XCOGBB9zT6yGvqqypDV8gczjw/3PhT1fVKDGRJ3kj27HCJjOOXoWVDKAiMFmRE93VaiYeTtDJ3iV
9rbqUkDfYZVNvXsvUU0Gl0LqP2PHlQoLooUOxJeYcfqkd6Ygb9QDufJBEJqf2NSRcDatKrMASHEK
reJyKQpU/C+lqkPrCRbz9pnxnMgg+ICfAPZlUeP8bFUs7TaVCUr/coHymZXltDmJVh7oncnm7I2O
MzNOZyRF6YFAV9iyo0acjJk41nUhModHxvrg5F4kOxbZW8WcCfuf/gr2XEJMFJVnv/X5IRgFtrxt
oPOjQGU1NmdDdCQIAN5yJhZqjr3f3LnnX7qoT5rUwS99KhHehqQ4esKGU1ZZanAD1aroCOoVGKZ0
Ppq7rM/v3ujd2uiXtUPTblrcN6DVPMhokwwP7dBPlMGKNOp4j+IWFed1Xc5vHjka0nAwrv7/7FVB
kBG+ybGCFrp9pSpcwBKWriLJYR+TgV58aySx1+dOjxctMnsuniTIQBO9PgKA3zuamaLF2ur4zKYx
kbzqo+jryPZ3Mj/tjOkPBqisvu2Rvsi95hvi8CnPnh2y1v+kwH8ZWwlVx8vTYn6QA3y+kgfiBGLr
i6y+RYqkV5w1euspESdv2cBYnpMC+QHbpNM4AotzzXxj0wbFzoeVrnWqeHXfHdpCzADLXIri62nb
A07ACaFPtJs+YKPdQW2G8zQwFR9ugSNgYZxWsFG7BszUt2UEdwgB/l7wqOu5EBf+VpwUec4f+MXi
VbkXDlU3ySyKgyUg9IMOvO+BB5XRJ84YvIU9OwcfB74W4BJZyXt+1TC4dZ5S+fCY7PILUs1zCAAR
XZrTSnoRm+5pm849WyFJdSd8x/sQkBcT2OLJ9sIw3S00HZvcHdd8rM17q8C6+cmXgDbVPdZliIPk
fuh9gsTLfxpnSf9bNVRpL+k5zf8MgSRpmx9Qoh3Vt38kUXVSGsORabx/xp7UnITDd8CSt5YBF3TO
gW3i+2O0ZNTh5/FkU3ky38Gu2drydQnWpijYMC7eONlupQrQG7Kb9aZhAWK7e8zHRQVgIa6Uk4nK
y4Mv/8x/HZiiWprk+KkqN/v8Du/EqCFLisPIUzvlUqpDJJLv6DwgSNpJOD2Vye3hEzgAjpP5sSdT
32m+b573H5uq+bAFq98TZGKdA9zZtHWPMM8uNhA5lbfDENpb/D3/mR0msEptoow7prac0q6vBwt5
r9ECgTt79PrvGYY+4hH/fOfRiChRKTc1OhKSs5s4u0O6ZkAuj+Tchsc2i+YL7TKglUxsS6r7NNss
o+z2jVmFpsSyjo0zKXcaJ4jbv2d3pHhrL77Z8yKLS920/+wdB+lXpSMIasC3WYkFJbc7FZEHJ2kA
uEKDrZtYIR56wBJ+oEUess0mkUGo8ZWIho67bKh6/RIs8EucdpWA61p/N/NeKhEBW8ZOv77EWJwc
RsbskgYvfSlqVvwSPq2G2nGRI2bfST9ACKpLuPlIFM3JNASTvRxdON2nfXCBQqe00Me7SbpyTTGb
H9f69cJeEnBB6DrPvSpGziCAuxbj6ikyogO8dc3Um/m2f4/TrfLNb/7klAUiwu65gmNpHiywxg0V
qi93xCjzHOPkwYCpjNsMmpJI5KybQEaMkL5bCbaWHEg17WGTXXcq+rn1i0B3MHDhbAluHVz5PzTn
tWbg+rKnHihbwo7o4bU3ecy+UnzGpdRvoGK71HLg8Wpwz/mx2KN9yfA/HzMO/qcwgVc3HPF8A2Ix
ZClIRVywLHSS+0fGyfPnkx1eCsyQvRkT2VvND24Job262tunCRIwI3hUhZSJbUUFM9ZdWgwca5cr
SkPU4qucaWVCXJkEQBlUvLdWODBNoVg7qX/w4Gy+W1QwKfNQJc6EbQgUu50FcRp0NjdoWPRtW2I0
QPkQeiM6aSTdHqPxhd9d+SDHoiluT6h2UqDWgHKdqrB6VUEY9FPDX9cOi7q/sWopkiCSj4gDMDZo
ZLuMQ8nNOovvH9+VH8k7jlv121KYe1MwO1tJt5GbnHGi9DgJ/fz88hE1YpBp2L9AtKBGC0HXlxmH
mS9QamoouwGHCxfQcHRKCm+tqtdF2OgO+E79rUlCL7gAJOUnZGK4756ur9yv2X0xIDI7Yq+x9OoX
hGS9qJ4GuzFzLF/scWXuCW532p63nd4pagZG8VqsKspn9n/oUxHfOJzYHUhg4cwoSlTK654vEgDf
imEiipVK2Agjq3ygko4D4Tdu9fyQZgtUftVBcWvuUkviO9p40Fom89E0hRrvwJpwzyKBmxhdcbm7
52DAyyUO68DQEzE2hF8MfTIDlg7kAggr1ITqvzF7RrTiGv2IQ9oo1Yc5xXV2STd5kIjEvk2ZeV7h
yPSw0mWjXqTmb7XIx9uT2Zzi9I0tF1awcYIxfj6bHoLY5ESW6jCiiCNDyhMRRpmSTpqQgeSnPMH5
ikoBBB7R8RWUuMMS/+251zsgF4eIcX43/VNLI6drcxqi9c7YRLXx0N9GYyqsVtsHts9/MLRcQjin
wd64CfqPYzmr5qjD2B4DRj8k3iOlUCR1dvzYoJYdgMR9T6cXLKPqMUQInjGCJfUYVrXVeuGEdTlv
mIgzsNALGVEspTirP4AMA4jXo2iDT01vm5JIL/nLid8Gci5V8OIawcqjG/8Dy0kpNcEnJdXhEWaH
fHG7C3kgXQ5ynsvXJRdYZYX1VNnKVQOCC70GpsXRMvWKWhOXmH+MRZFSQoLgtTBAeiDCOHaXajz0
cCYUjD2yezAzySyqiwD+r20Vb8xPbCOzxudmHLaBQqKQj6B143JPloQeQo/2Ee3TMRz3gG922biX
k7rEmvQDmGZoCe8dTmeQCaLqUAbDyHTuCcG+kEtBJknJMju/RZz6OrCfYld04gC85xZ9oozz67A+
JGKEwjW8+P4wftgZbqL3QbMB7oNz2/e/jnEHY4t+9BEi1AygXNk+pN6CsSfI61XzkHhsA/OA2OTS
TAxo5DHv+WoFK7PUgA08xD6BSbrlUn+FSHszfPZS/w388ayN0QOpg5qX4I6A0Lu2KSdjgvmmDfTH
OTD645MQTrwpkRvVUh3d6F241WRgITAQ4syRSl3jfdcP8NT5q2baYPnambnOPGaV8KeHwhKrYAAY
UfY4jOk9RF18Ccup6OAqWDELqVN4Xp/OS9LWDhPjP8Hcc6kgmQ7uGehNpPtZMyLdpd4ED7LSTftq
8hIdYDwJVr9e4uGz3RYZUeGqqud0ArecnbKGQiPL6TkjXd3Yn7BN/dyKy91kvCzoz2NpQP3EjGff
U7hp/36h5E9OSCXw/YxCfdOAj4Zt4RUY4er3YC4vwbGp3ZMbktuTgclo+9ViIpI3Qfo1DfaB210w
Jly3lm23U0+dXrAmzoTirCmhz6Ds2uXFC6ykqh6bPtB0pzwjQ/NLXQWfxvTBjVqO4vPHAS8bkx11
h9ZHpxgVMwLGht3IGBgpWzPlm9QqidsORcXCi2aC8NSxkZr2636WY+1ALcMui+3D+BjfT1oTXMFJ
PWojR52xF667CJHD2LzSAinbKqZmVlUEKdszy5G7jGdD1aA3i9re4gj6e+/7zsG2sEbWTfp5f5Tk
qgxdQ6F3dczw4p7VDYP8SLVXDC7n2kDcf9DcYcAyxL6kMdcKIBJE3dKijRUGVIfOdSH7pZVF+gl6
MqtDas8VYtj8hQfQ6Q07xQARRIVZe4YjObjnMinR+Je/U9+7etrRwfWAMIFIL/pAF44/iN5kvrHo
VhXfaMrRopAqev86kGA5bSeFVV0BOw5Poyer9rjmFBVXswj7jYl9JImudSjn60USty8U6P2lyb1C
74vQVct31QdaiLI+By66PYi0kEox/pN97DNosmtLR2h/fahKZk7iJhhQ+lyDxhGGnvSg7ioXIHCp
BylO3g2rIXBmGQhTaSJfXwq4oscs+syjy5Rh7ZD9L1UBbcdjPn3zhN/M337gRpP8aFQfGMvA+3e9
vAp/XtMl3ks5yOPXs4Q9m+vfGCfn6BfWIy8MtcWbD1YiUS2s0W0VJDx4el3/iw0V33+R5q9FRM9D
rdPhOBS1MLu0Tunct6VG/zJ4B4sD4QCAP7iGXslStjZTuURflR/EBsxdsXyCJf+jFDZKKHWDKqbd
VIqqAIluDX99nn7qfNpcPUhOdwtNNvjPtfJU/FJvyTmy96KO0bIIovjsZU5UKDl9/6lOTAWHw3cv
/X0nglSoksrXa7MH1a4M1mP1eWq/JP3WKQnpmzys6tuzs8RUGg9gRd0tQVarOPbjbzSw9vwn6snl
UG9T6pEo2FBUHxq86IttRTbwwSvlyxkzedUCHrMIhfZJ8eW2Wdl4MQ3V5JELEHJBGWhaq/f5yrH1
kr9gJG6X2UXqzIlwAib8stUF4HcD6eJZENrVkv3fjLfSObz+iVqPBBo+SHridJ0mAB0M2LwID+RS
dYZFaNW0oj60tpiHFp6LTYZ4hqmkPbMLdCQayIWqnsIKDYzYckvqf0gHzUTTUp19RYY2xUjVkFt/
gS2atyi6GhZm019lE2hagDWo6uKd5eTsGk2S+y5wuIJZhgFgV08oMkRusJO4yPmSjO3hAvCCbn90
HmJklzPDwDmkZbkbM1+Un7D3aeTm7hR7JTdF8XxeWepfLFFp37qXPx1pc9TYk+DX9nrID5+hSXB8
h4m7VUyB9qyLw/B3lrEqwxm3h7FUebd32b7qoRfBOC+69j0sA7k8A4Dar67Q0bER6ugo439XGr5N
ajiNwd5Db8ERLzZRIpO8qvD85EaalOwHoZM5SrIaDxwX5kbXR8SzpxnRMDOkSP5hJ5r9/DGmKYVp
JmsRgnq9eDm65PReQMNXL+UAHg87tIsbz4Iy9Y517VE1htyFW0/UP6PHbVxLXr2v15og3sIpe6+7
55qpkpUQAFnbNL1PIwWkXsLqeW8CzL5FZhbvo5Cz3nxs9i2WHqJmXKESEyAD6aUzU2Ff8ydESI6M
5p3eB8QHH90+jTo9JHeHOzTRUqN6k0hYxiidyKxLRmBLA9BLG1CklpURkU2iLUumGV/hdo3uCB3z
XI8YSfPn3DfEvLmlqkY/vhp8Bp33DrZtmUFM5FLnUKTfsXcW//0QFP+a2NpR0LEWKb7iWy1uu7Tf
WHiFeBkF1VvOsx7VA0NcqIOdO0nF50v6Zi2hCxCIIOd87QHGgJh9nmYZUfdDxZAmS4WdNgnQ7r9o
nPBZIHVpaPiBZtA1S3th/BfXqAoReLuQKNkItZo2yHLbCagLkEp09Q1FVn8nHTmdnHXOXkkYnc1x
trUyZEVQjVy6fVhjf0JCr/jDJ9puoQkFtbfySoQOxeJh5P+ftEmEHKQKs0k+l+NkimZAeVB9/StD
opLQm3NwlkBTVApaDWaLWFCNdXi7Dbd5qTVuGv+5IAenmGkz8DDz63H2h4tUlqg0+x6gMHgXTYad
CQaLEHdhmbCppl5CyllzzMgeIFGG5ShwHLaWi9s1MzHPBWTDNAtP6dFtjuxg5L4CKT0Q/BJuawW6
MEhotZBYz3883KohBzwsXSnZgcXqzNi9nTcLraMmJFuLxataXfEkHOSNuXEPjQiv+ZeYlGN9sRlg
BzXhqeyLRUhAvJDc2buUylKyo8tg+1ZAj/G+HBaxFfGrE73OHl+2wL130PAICGWTuyfu1xncGTVT
j4TkRkCqs7LVrVtf3NvXWYX4r+pg1np/Fa3rT4rRnnr1JuoJiE4Kt5Zok2m3Mhm92F2jhoR8X2es
y4Cd3c0AlzYd/hRrSoUhTeVJl1m+In0HqF78ci+x6b9jCnVWuvr4lKD2ugFBkg8qZPUrdoEL1gLW
N4Q54maVjT/TmnLjK2rBGhMdPIpcGMbLRE85UlGM2QlF2+Zq6btuyJ21aWvvjIXXgVT1xGtGfvmW
SmYxGry++IdM6Le0g+76QB+kuXffzLSeY5r9/Phg6n5NNsNrf+0lzCeT8mySNq9530afpCKG9u6I
h/PR1iY2vMprPQCI3fQylZHTxWmfafVrlwDGFfl9D8DnEbIs9uLINKXpARhJK7zC3eLcjyn9UY//
ab7lARRZP9TeAQjJuoMcKVy9BzmxpUzQgRwm63ElSDz2Idt0/sJdZEGs6wOX1rytaV+6mhDei2n0
DCWs1TJGIEogt6/D7ReSkOntOwlZIOZ9RBaXqyBQEFU5Hf+zRNOmfbR3KVem1DABXPDMLRoGDcWa
yY06mXhrwDsfPP14Tugu3PpOgaP034SbnvjB6unxSC3AhVhxD/tUWSDBuCXQjPZ27ASo3R7ezdmU
PkAUJ0RKmnlnK8IfrLlkLC7CmDFulaHF55qbQME0AAkmugdBP2wxhBCmoSiVgRrIPUIy753i8APv
VHoOGQ94BQO9B8DtgACrOajREqnRRImZdmmNQD+2Dy5rCLF0x8nuEK2miBcSCwA5x2rtejUl30NE
Ab9nij+tttteO0U1sXsewm8QNFEcdjEnrSAF2RNRDtK32Wj45rQpEcV6Ff0BK3bKj3vWxUGDroIO
PW4URASH0uMhikj4xPoVqEuw4nLBbcXjDBoDW7k69f9SaZCkcfKFBeGzJeSatDX2kBZOYSQyUVDW
qD83Yjmgv3IMazWlUk14ZJfCM/RqDY38ef1RvXpicW3vr01JyYmOwzmUhQHkTTGFVCWOhggaC/4o
M5s786Tqy8CHxx5k/jHIouIVRv0mMDwIrIqX7z7J9LW9qdS3HX0OuNRrL/4ZKvqbu0+WABGCNv6C
vbpedxb095erdKsdIb21hDie0bGbR+OOqsX5Sk6Dte2DWNl/+UR8zdl9ExmgjrV2ZUlDiSd+9/BL
xgU7x1dEnEnogeHZH9icmyLsP3wSg9e3kIQpi+/i+tUAtVfgVGlwZT64PDe0BPWgp97G6asmYPLZ
+PBLd/q3MnWR8niUZrNA0W82hSvSzbGqxfRgLgiM2PTAcGEBffwa3W2p0eLVkDLGujxf2K6KqDQh
UGicChh3v0o5Bu5OXrSTZTuryxiOC66CSDV/snmF/rdH7EoqwHAKuAuyWETxM3769fZBU5pkGrcw
ImKHYD4dPM51bxkE3M9zuWF1gkT3PFoaXeat9no7mFcX0+V2lT0P3k+BZji1TCmNc/ba+evubwz1
O64vF+h13o1H5AWin/PgMToogOaL5XcAQ8x8F0mF9ekSRW9db2FAMLHKKTyDvG3ODcWedKYbskun
zfXqZXYhXS7T5XsTp6dy34uu+FtaueXMxO3U2AdDuEF0YJnyiFarnzz3ljOAmEgsBtbUPRSuXCQe
/x5LLenoAoKFvV/jOvx5Hl7N6nmtkkyipjUdnMVLXws6IcaoYPFrsSX8/zGzEnhM9X6PPfamLS2C
yFnhNQZ0ZULSBTp+lXxIdmsU/hyRDUh7EU93tg/864IwsmV4ZigSaujcaZsvk8PN12rr2Z5USdVn
EW/6hBvMIvsxdZeY6s28JkWCFvwlT4dHxihg+Ygywh6Q2iHAxn/emvaX4yhlEHvtJv7dAnjCPQ4J
RuSc6FfGeyshVIFX1Gx3LzTKXGs5hqd6jjqVf6frNY1EV9MJpoW17niiqaB8rZmitjEOW4ESUbpp
GyXBqUuyW084GLs6w8it2VZIbGtsnMjSqO7ccx3pMhc3uZkC+vZEnvOt+sBGd1BE3R5y2sE1CIPI
VxgKbOwr7w6L6RtEy5vx/hWUDAykvKguFUQIG5g+MtN2vcqdGTV9FzJsiKl+VgGsdJOUv8TRvqmw
uBt+bIW3h7ijzbCjr044m+pvpuJyT8sSo2PZDqUILzw5cWsOzUYNuYwCKXwDSx45/Q00Km3jA6/d
hyGp/CRtU2RwbLFZaSRmMAFV0JTj6hzAG824YyxUNnjn6fmQk5QuFarmFn2hYBytzdklP18uY7UC
Bp7onleQXsoQDQtcKRCVOgO1WmX4pO+Ii4NKe8Pz4/qlDmwVGg8OhJGM3BO6u/n6Pjt7Zq5S1rdM
ZG0AiBza25PQ9XEMaZO+HT/QkmSSQOhGCcAea66NXyLR5MlZp2yzz3LZbrMkq794dwHb/7LJWbHw
hjPO47r1sUF5fkNM60NdXo1Ht1N2N2Jl4NerngAVnJkRyDYAcaaBu3TalWq+fcpsKOfQNHktxyCf
TQ+R3DYn/plLpqCUtmqXoKaTnPEGiCAmym1wQxBszf0buOEGEUYuxnc3LlnHoxUmmo5jJAbSll04
JrKrQSNuJpUp8Yy+Hxp+xrH0UhdBVWeU1bvvwoNu01x7ncD8xKEgz00QQSPethjYcfXtVm4XcsuW
/1vlnK+u28lL1iULZdlQiTc/JWIjHwnto0nJItEP82+uclyt5qbctZkoUtsVUfZs/UL50GIS8T8t
2NOfoQ9zJ2HW6tuwBYjrPUAxJC98IUZih4nk4WTUuVQ3JDSMDHSjTpMxyzzS9i4cX6gbn1gSpnxd
fY9UxOT9+tFs2AScFWM0Sxo6ZAN/I7A/1WcJqZB1mo3/vTvWRTbaldRAk8hmVjok7w2jh51Zah5u
Oi+2JTOYl5sO//B21nEMQQRQ/HFO03zVTTdCnsdOZVBJWJ2UQ2Vw7CqC78o2qJjIqb5zlhk0zPD9
KftateoX17XFO+wbCT17PKXRmqOGVcvLrPHZNlOpTc/cX7Fxp9MLa7s/4WxzXq4nypQ5cKxgsGAZ
jR5Pk+jmUGiZy25eragqCK4N68H5Z+pC2JF9xcSc5ul/OZJmALIQ7wAH2PHFuvoahHFsaIZwC+M4
E/Hhjrg14tuf6aQCguFKBNyR6kFjtx7s1KVDCvKUdAYRD8E+in0P6zygvQclJwPN7Nqt85ISrIPu
ZB5jXEdV/8jJzEILSw5fHkzS8zGJYm2IHEsn3jfVZErG+2ZKcyWHqoaBo/3lxYPpO+TZP/jqkGog
xBGOF1kOSue7gtPb/nTdg4Ew/tAHtrkC3ElxFFWBwp+MsSzA7wgP9WirhVoq2ZBH6Xowo2LrHqCR
1r8uTtqUbYxUoVM6goEZeJeog0EMXoUFSBIcr972YKsVqB/Ve3DrNDbXbhyS5QQCTqeGA+cEkZi4
vjGeTKJf1LlAdz3mkiT5F2NUHg8eg90UYsZleSYhzo/Nhod63NRQ4KWucZSEb+s9mGyrThCqMPVV
p4axAEP73bQby7nem3ycgIZTzuefG/EAo0p1pxnudhhfG4m156RFGcKtCedFfsGf4MOs5a1UQnqi
+/7d8Dd/zJlSS+ChkBWDM3pkKjGHJUxh78uijXnjTlQm9Mr35AQ2hsioqLxA6/2oHvOp1OOXfo9t
AJtEyr/vNAcOBpSfW6wrzQR7JKlF5V6u7WfppIqiKE7FMOKAH0ftI6wKNOkVMjAATOasLkYlUT+z
t3OUXTvmO6oYYhy0zu+FJmuqJa43RoVtBGo/viUSenkXa32+QmfyiQeHR6+KNuwlgzwQ0WJEwzo1
5+kJL419BF6S0hBSYnCYom+lw1fXm0FkGd6Ss+rqihJ4vdJFeeEjnt7DeNgoxEfDgOHlU9SbTYX4
MNxWHJQsMwAXZDeJmiG7qlq00PgwbO5QQZCXNQvCg1MFPr8SoaG9bH5p7UoIzTCjpdmoHS/wTVoT
kNWqGLLU47KNoyvktDyIr7HlKNQ29QHR92sQ84YfySwjG/N+bH+cC67GkGq/L4SBKz/Jnv6LTD6X
I4O0dWFIG6L6yGkkrCD36kCkJrGMoOUSTekulHWP9SYjZLWcKBK7jBISSNAoGaniaFA0lUayCtC6
XHykBxfsV9N/ZZ/iYn4b3yyGHb5UZfLX2Ik+J/33IJRsWzpkJSg0Ildo0fttj2ulFWRDKtJcD5NS
naPF126cZoju1xg9jeYjlVJhjl67WO4RI3aPk/uFiWDhLg/+wK4X0ygWZcVW+x6owTxOKDs2mM3I
TrfPKcSE+UzMR34uArpCGpdGPf63dXF7qfQl7i26XVhTy/vhAzHaaifC3L9oHIUBlp5A9pnvlScs
ugPqiY5SF/KA7QQtvx/sqT9zG5KdWqwqMzRyG6oB8iV4a2Mla6OnoPZqBvFTxkK/uhBlRh0QKNVz
IcccZArQv0Y7dKyMAQG+xW5+oEXB5xKeJGu7GCylCvsSbu2N30gkqJZcfjz0mBVM2AXQzcXGINlC
wEoQ6n2vJyJHkX0nIcnCX/J8wi+t3TGg7mYrNPcAvXkrsL9vHzanF9Y+e17bGu5Fp9gpQtFRZpws
yFMKhl9rPXqByTdv5xJsjpKI+yrC8zwVKQwjaVGfShuSwhbIQnAzyzJpVZdBwKEBFisBZhcvovh+
sdc+FhwKh3ldaGRoGeEadnnRhbEhFc9yRFVRCyRE6bKweWlfRGhd7Gtei1e0aw8+o0Iy2Zn+jKo+
w10/Nwcl37et85P2tmff1IFc7TRsEzEtzJvrctsC/pUCqBiXkHusRs5IIZI/rtzaZnvtaikBZUwY
yVTDWjiSi0192F3O+UOp8hrMntvf5hci7vLafkf8ecU2x83Pmnpy3QrtAD1ZgMb6FviXa3gFOnH/
oep4XUXUlgJ8p3b7PzG8pc4E56VThgcS8HHCpfifWVR32aBuzDH3bdtbMSiLdz27oVI3r/OKIKUK
gIgLtczyY0B9Yd/PU5pWEhETeFXXUNaXkinFSc9B4LsxZ0J2SB75LXKxgyNXc5sLtAk3SFavRd0R
LvKIxdYbFuG7TcWBS3Ib9A4Kky+FmoY1buyAg4wjZfVLkYw2T+BG0GAlzNGtDEn8zifNmKfVJmfo
QHFOnfURJInsd+1LZgUwWscxEYUZHP0cLYXMDG9XsbvspCbHe69T1Dce8HVCd977R64zlaf4NRhn
qAy0y7OmE6q8ZgxvkMS86r/3mwzrYBX+lCMltsXE6jK/QW9O0dbIhG6WSRgqI0NNeF6R54t+7YMN
Q5MzFZv8RdiYx7e8gbdoztEjHzt1VwSsPRHz/yZ2HgnPVRPLn36p5aw9d+aPpuKLues0Bya7OQVy
yRKoCl+FTXHZHOrCCMl6ir8gmOCA4/p/MsYkv9VzkMTS7v6Qm6wXCu3ZOSB9/nFDwJkVoq7LN3XJ
Ic/50Uy8K1G96egiJJ7186VvLwbP0V5I3NtLb9syXsooFSCmIPNemU3ZKJJDyXyzSRiEl3Cj61ls
ZwFCTUSCLSmrdcTWdWR15u3BSLmvQuew2edGpy4U3giFfp5EP4P/Trz7cL45eWN9zin+tl0qFFA/
ZrpGJohxCQ8C8PUNiZhmfiv955ohLPU112klxmLRRBe0V6CLjMr1bzJK9kbrjzM+pUd+jR/4vf3j
ANGlfyZ6jEmUmIh9dqtSrl3LOrbxTw/PciQHaaOr/EWg1VCb7oAxv3AesXbruMnX8PgvmWNgXn4c
vUsa19c6p1A9/5oXNU5AT59pKM1LA10kXVRzgVkaYnHF446nSB030De1fZigXO3sPxXidNAup/mx
FfFoMBckhOMiiInMfwnf0HaFiLDflNUt/9+I00KX+Pc+bw8FUTjUWvxtTg9oQu84ENJ0CnUFXLyQ
AyzwiFtQdIPYGSYiEdITGrpkGjf8I1K9Y7wfIUe1tiimcFu6baY6nwYGGd01DCJU7MIuJBesI5S1
AsnQz/KfFJT+k6K8LiNzEiUIW5QT5c6pnsmmCPbU0oj0hTJ44V5kiSmEobsz3x5/S9EBWVbZ3X1y
M8sx5L8DQLASIVMn92gVq/CbcymP51Ltov8Wz0TfxNiSvV5WEu5mg6ZltVW3s9kdG0QaAFadBiHj
uAf0Jit0ujo7EbN9YLGlzkNjLKXsxlfe4SOuQ2VwgeBnFytfM62QxsQR9Su4OVzwdb17/vviFyG/
Rmu+mJ9au3+jZ8Knvy+K0ccW5poqca2HC/jPpiElswLbgyR3o3fiPj4SnFDiMgiQopJ3amcOKRbQ
m/eY1LuK9zfUP6unG94gi7gA6K3w+aRZhvChgElyhFS7mjXk0Zg+oFwx3+djG1aF3bbVsqK4zxG4
5n/0yjuiC/q1YaTGdEluBwkH6Qt1kdSy2EB0+KIYCE+X/gcdqDboSYjiI1oooQGSO9YUUCcV4GEB
KOKs/VoOaREr4k+dFMSjwbe1k2cCyr5GyrIzKOonoOYE3EiiLhe3oeT+iia7Jbn7WoY8xlg4jbps
+Tvj+FX5zoKrgxaGQfAE0YwtS2HEyz4Oeno0nlBlbnJtztepeywC8JoaTCdDh+sWOdUFzfyRtblL
m6kwvDJtYkKeQGUl8aulSKU/empsdO/iBUrhNRLeZAN0w9IWTm30X47iHdP/FqHL3pAB6icqnSHY
n26TTR6sDy0qp/xXmCF2m9xbrxB3eAUjW+GzLHVeJE4gB0ow59h9DdjHV6paPDVu94KB2cCaSJU4
J4+88WTKoM+ZuitQ0DqPTdbgpw1L6sMfnRMzVWnCZ2WsxyJuQMwBu5EBge3RNpElTAtbOKSNaG7i
BpR70aqJnYBp3SPZBZB3IJBHF2FOEXbTJdYuCXKz8M74DAsophDfryW5wQ8HPnbtvIRDCXeut//C
WWepnUKY2bBWhxF2Zh98pgkQVh9j6c8yhcQqWA9UpfCxgpOix12Iyi6Vkh3IhORtyfMquNIuMDcR
gaQmwXLndJnQubvliH1KEydJUaPKJTe3t9ToygNIWjhQkVZ5mHWtRCtrOue1xI7+LloT5BTvG/Tb
ZCiac9Ij09TWtpuKqj7VjrvxM4JQslNhvwlHDZI7/GardFFF8v5iJPvypQhmMzzlQBc/bbYakG22
xmAI77zjN/K0li7rqmrOs9Vsa+dSAj/+Foz2NDpuaZP24W8GD4TRJ+rh2ycbk47x84ibw6Q9qP+x
T2OxpAg9QUnDi9hjRlduXD3hXufnHruNmpxnDtHdEO31mu4tgnKO5s3Cym0e+zFp7L4C56+Xazcf
NRL1Fyn1Hq6BGI1z1v+iC126/psqeOP3lxO6Uq8uS2vLVt8gnToKU96w5yMO96obindrmu0cSM5W
iyUrbEyfbryX7jTSwTCmpSzOhGW5GfRQcruq0fs6O7rPCarhHHQfUraCSw2gW2fFwuLfe+eFDg14
8LKyMmTygW3X3Kep9CguBwu69fL0G9A5guCm2DHrnLP16dnL437T3Hd92gePhgo2saAHRtqW5MT/
etrCvIcfu3us4t8PSGfDvoiR+jyuxh6JYAKNbqBHYUf7Fjrq08bo2l+QE7CSwJrjditzQq3FQzDs
arRjj/plXj+/d/W2jiEc+xaRAwj7TLXjTGHB4BEV8X9jATwxqU7+Sui9I+cQp5VQw7bmOp004rWh
FEk/R/6XBZ5qrS+LJPLks/o3C13jcQYbtOnyo7q97YhHpBBLr54ohvZe5voer739Sm15MUxlnQ7c
XBWsVTQnRzdJ8M1sFvhaJymMGZD2ACHdsfInoPBBaFFCl+z2ZE3vRqlMV26SdDt07iIKWll2QYFW
b7HKK8QDK3iRxrMA1LAK7lzGu1KI+Mz+GBmfhpgQ2H1loelj6RualLW8/FPjgKi3uK6H/+E3i15J
ASsjpN2dmlY8kV0tZHiX4dSycTaOmozncASSyl/C3b82ov7JpN9FboMX21PJn/K3M5zoyualKO+h
XYByh5D5Ii7yUfpbaCYOiGsKdjndqabcARfKj/mupPnumFGqnofUQCOIDcnVrgLcGRb+C4hd6mrP
eDj95XSP2u181gnPGzVx0BH1IYcowKQrK2It4wmfNJUlNGE4B8L9lXJyFcz3vUDI7T1I4I9D9ZQY
BjniBc4OyEyOf3JQ3hB6GW9If8HGPifu65ulfWrN0nxLtvRqT7m9UtsxmbORQt9V6xw1YfZjO8JO
G+krxwLuV4cyTPl1dOsgWcyTOR2OqdSnxjRAwJI7YZV4Egil7hK6ANPQjXMu/5QLszobUrvmule8
kvgNUH/fdTWs5Dv35DARDtPjU4LQAkgtOqquNIya6sTnF6gCut6tI+QAsrx+zj9BLY0SVGCAY+sq
VfGQFxT7CQbPr6FsqnKYXAQe4+7ZBMGqzZr/yWXTZ5Q7IJJClzAtbf/1LFrRg02cKbWN1wlbEASe
nYKm1GasIPr2h3fH0f1GVRBP0etRN1ujawgj5jsZrfG+O7i/MCJVRamh359As6wadRacnw5ijsCw
PKmghBc441taUW22yoC88A85ZjdySq92LHsvX0f397gsvuw2QBDLeBN9GY3L+GeuX6gP0bt+GQkb
tA5e4GMQE4+hf/O502JsbSBWDUulHMZS4uW3/Oln2qd/39ivMFyzuGu7/bO1UtbTCSZ7/lP47r9p
9W+3QVP3BNoLcfsqBxA0d6r2+1614+PXK1mjQiA1m0Xk7pGVrvQeEtwg8V48YoQCLkUiB2qFfuXf
2pVxypxF/N3MnRLzxpRodUlL9BZRmfN9FmyqV2CfwU5G0uHTgeaIu6M/wUxpyKDgVm+CL+XuEpcc
FpoNuIdyLkhOHk5XWRZfLtDT7GSS9YvWQp0E2VwayL9dLKmUy9a7csKZlDMihMmzXW/0DNC6Ry1g
mNdGb29gcSwdkgUcDEi6jRDhOWXIsLfYgptptuEURd4G3RHhQQr6DLMhQVsDp6OKdLphbHBxylGW
IAz/CETlWKnYB7QR/PUe1yjePc5mLlO8p6q8nK1LW4vjCfsNf50hCYiLE13yjzBQQ7n8I0Dhw6Tr
lJy6rg2xWJCcooYsPOtcRrnUwv9sPCCnEMS/nHrAZhUlXtG+QNrRTyz8AIPx8zp4Cw0NGyVOXZCJ
HPvGBKv1lG9cH4nfTRC28fG8tdI4tC3Kyw9HfNp0aafCDCE661Pqp7XSg8hQD2/QrnO1cd1LLkL2
uVc9GIB5BZkQ/vUeaHkHpes+QB7G8LzM9zPZzMljaz+7At3UITgG2rYtZfCm68VmmnYy0/c0Ts5k
cILqRwY+Dgne33HfMSq12rOB+BMUR5mo6OwHu1svfQ28jW73apa8Xsfqlc8uCf41Wc+rzXFzUk2Q
y9MhV9VSL1Hp2fQdZSy+eBQU9qmpwLcbuc3hQGee9Pi5CFHWcrY08hLySMMmD1Myz+RVoLfk88Xq
QQLNf6nTDG98X2BFDm4Mr2p9Q3a9RAsgmJMCzWAxLTvQDWW2bCjseswT+PFDJRcmRixihuANXW5u
vlCwKPc1NOcwOYxJqL63bdVHya/sedMnTykBqsJDt8XVOKKIml9+q6VcvS46MFj2lzgmMMBxsplu
cYm7ZMP2qA3AYlMOF6Smcz/aVAhwxV9sY1jWzOW0wTknw2j/qEjiw9tDmaJaYBcvMHm9UdrWIQlp
eCMDcAWFXPhoW1Rp4B2wag65tLSat+Vye8o9fHr5m/jhA9Qxntvx/8DYAI+ZcPLzrc8/PQUtfBxX
52Oslt2zuzfQaNg2Q2h8EHRwlINmglheDUKnhUDFkmfYgEGEbI2LMD0tb2tD12j7atkdeDJOgh0s
UVLm3S8+FbL6qdpX/tZ7/3nArdiluVFqusuTxKL9fmki6XHntOldSJ6UAKjx7Cv9sgRyzWhfJeg2
+fC/ef1EtzCc9Datdam6uqu49lW1Wyvy3+8WGloMSeH7wEdsgP0XRBMb3TlTeUYkVThjHTa8+5MI
xBwQ00WHORC4tYdxQ0YAFC9UbVEm2+Y3AG9VxMaHArp5i/Co4VBrAkJPGuq/3U7g9iaWp8+1RoRj
iST0D+EMsUvlXzTWVpXkG3WZqGPKKzghMM5OzVMCqHQMSc8aDLh5MRaSQkpTRsqse7aANQqg9nvG
72QbByUdy9eMOKjiYQ7X22VMgCVtzA1ajxzbhg9Tr3RaD8Hxmfqlkr9Y3VsaVBgWh4w1Y7rwbIBI
9URsVjQVDV/KjM9qFNBSIR3m9rSMkXik5DU9mv/KDdkx61hHhWfwDOARozY9NcttfurVzafLyNWn
8CyU7ONxYVVz9yGYwDwVEfpcgQstDV0UmFgfOc87kZ77Lx4Ul4IQ8q+7/A3YGxBg3rB7mbhIFvSp
LtP4mZbQ3a2X6NFS4sPR2qnIAe4YXewJdcOrOKKyLMjwPBxTG07urXCc6a7E3QbVteBQJSBnNW60
D5xsBoVADrB1663DLYyv9Xo2UA8xn1TDNSZQC8WBwg3WUKWZqRJLuFz8XFCpodi5WH68kkOgVs20
zxEdSSyxzpwIYRMEmeOUpKKxn/WIxjdzNbzPvA0tXS8Eqphhi56E4s5hbLMLnTGUM41a+Y+KGdn3
6aU2jzwDFB+4GZcMZtKFW4aUc/z5Hyqf7zDX6jU/RNp6jT+T1l1xkGIz+BJseHFgULelML68Hy4N
YExNBCjvbasNW2KBcyyrRqxU4/8m7S7CWnUyop6xAY4O7xUFj1v41FnDFiNBhL2021Zy9F/7SJ04
LtpMKLmtNBa5QZMc+3ztGnTytxfe0Rtc3Jc4ceAuvSgCAiADlxaBEGiZAQAfhsyI8B457sebZphy
4NG6JRwV8aWUpu+mqdXA2BmHDg+yqrPnbNC2RZTTk9DyRUZ2GEBDDF3Rz8+dxJDn8MD/4xibXkgD
s8YX9wO7GCUrRgxE+MbmUi/9yYJAv9prlJNuKUzVt4ZpJQmD/oN0Sc9ZalpjyyYPRSUvdUzWDndp
OnUt0QkSvk9j1vSO5cmfFRdu/spOMMMFiP4qJ7PmZrzF2Bgjb5ehAXvNsRknhQ8iSM35mT22ibCq
PAgUEVrjSfLZ/JgR0zsR+RYrkiacTFKBAsmWoC3E/d/TrNxXBDmYXEVO0rqI08WSACYikATAETmY
9xX4rDdh8T5CvkNZYBBPJ7Oa1gPCQx90mivAk3Cvpxj2s6sF2gI+9aVhTL3NwzXOENqIyd1dcTwe
ywSXNvQD5X5wLYc4riYDHCvvvRaRxXamfvhZGx4QqfbgI/H6UEtn10gowZYYMnbl5F3/Ki6qg5qk
8OvXWKr+R9s3zlg/L8YiPnm2IqClAaWtXBFzidgB30BYs/cBz7+t++OiKSFSGy1Qr2gHElVCUBLN
2oqOl8TX22y5Ly8CtTfYMTu6LujpT/Aq27m11m5hO4byav/wqNtRPGGSL7TEDok7+7uk9fXieTlD
La7x8roU2MrGQrNd+vdWPyrcVgZDCThziZyfgVWqZfidbghcGhz6LVf4Np0d5xBdLFUZ0isH9EBO
2/0SKy9mUPIXNcwP82G4KGISht8ZVBVdFR9xD36tt24CoqEieeQLNzmKbUq8E4ZFoDjK8Kns9w2V
MDGwQtQHnkz2OXmAGKsJpJ4boKqvVOHw4gYvzcbddrsbQmq7Z6iKjCSGYMvScLkUqjgD/Es9vnxm
o57WNbtihT2qMI7ypPyFsxSj2QJ303egxLFyQo9ITxBE0KS0ymBAmiWae0GjnZcgx9d9N1cMzt5f
jLBgd/lgoD7T1UpJspFrVBDpaFjM1DpSHecoGs5i30yooLIgZzPVgj+QFZNGs/OJTMppT+93HNaQ
oHjrKAmTcVNP/0elS5t/f+9af9Obz+iKrUn1SZG8tq73b45+m5lvYKXKH1c6Vk2ARp3qRZQlMotk
NUenf618WqgQMPioLzGfmRkZGQo9BB8pg+8vPbYCk3OunWLwKU50jBs6Vd3vR7L6ajZ9x4CA84Gy
4iGovp71p/il8oBzb/JT55LDme7WnIotXXSpHRlvIzt5bE9XlEeGmEzB1uvLTdM7LXaVBZPZnVE3
jDn01H0RVYeS65iXp5RB4DRt7j7Uc3TBBXuiFXMD3NXum1y50fr1mc1bIsFQoLHHwDBN8qNFKy8w
PGqiJ3kOfDNTTYSZWF3ZNRik8GMptEU9Zfqjtw1wLjMPIgCyIMEL94zJ3087cv7o6q/drA8CDL0Y
wiM0qudO/S2cxrP/jOQvvhGKxJqAj0HcK0DouU9Fqlzj22l3z/a6QSi5xGTT4nquCPyZDjcNduI7
Nk5k+X9QZiKjRX4ruHwrhvO9ASPsQ/uJ9ItFzjWYOwt6rzFF2+pj7xmLqOxbe68Atg8LetuJdHHu
TKlq7dj/OyBy8B67czO0MUPWshon8H9ZWwmgfMitMw/2wsh62scs/9Fx8FFzV0g/UitGB8BOdHzw
rj+DYD047y2lW7kMxKIObfjpURdZ29941qiVxCI7ySwfIEgrQ8WxtRA1fU5fKdwLmuSotYL0jRFu
LzRt3V28ZKKg2Nau6Ayz72rx3nIz66+Z3l9dKeizj/cJI4oF0hUqr9LlpCRFqm8rkRJPd7t8Dnsu
Gy1Uwfvo0F8HPGnvHHqNC3XtzO4HImrk+L+FFX0rwPhyQu558znylWTfLSSqmtm0S8MRvggHJCaw
zJc3RC1JE8YnmCz59r3AdA0PDY7OQsCLJX1vFEdeqUtRskMqYkjKilgBk5lgHuyh157ozxWrYpqk
U+zJ0e/3tWQ7o/ecezl1OYGDbp5UhS/LUAsFp48oUvVxLDlOnWC1GRDYTC6be9Txn5smOE/w08f0
AX8mI/kX5P5Qif4sznbl5SIFdhWHaTIfjLakwvWPfkis72ZFv8rFt7MbI4dGkhl2FhHrA2growpa
Jqct1rLcbcV0Ij1B62PHAv948u3uPf6iZPqJQgIH+JFhtZ7pNQC3GoX7mPedWtSNR5+jXw4dDYHT
FRPg5iFi3mAfdo054WUOGwUuni7gCWY67ZRKvjkhlu1NhDJmNLLRddB0MlALRJKjZk9b4Rwjzxcd
1CTSfkzwqT4xi/409zMwFMYapjDJzxmzK5tXCQZ6qnD1nKnXIH9wPWGuur7GG+PcKL8Ui+BDzLBD
zd37j4E9qZfRsugjJNSfVqAxebgrQXRQFK0OgzBEQUeZBfmqgYQUm/ogpaCVgYhEwRgRpfbv6wgz
PdENvASJS0xJHNnEpguU82Bs0WHcu5HKMsdXFfS4juisauDUJEdr2nXd4LDqZOi82olADkrPgXbl
WrHyYF4OiJG9zGyNXJWx4io0rTD9GC6DI5YaP1XpeF+Guo8HEX41f2zXIjYKO304pBwZo71qmxfv
mqNxbWUnvXoGzYcyiGmTqDklBeT2xxKFhsczZwtkvM6ckQzJ7mp8TmvcqeK42cbA7/i3x6qAtqNN
UmhToXMlhchIXzRsFsDYTghEDSWEmXV/0kUIPeB87dC7tq5owOla/xQLLOsV9WQc54Pem07Cdn0G
iwTT4MxPEsuwffOR5vJAGzk152abIfA8VE7HwecAjKiJLLSczxLh6A9ybGTaoKHs2e57XkcQi4M3
0Roas9vj9SLF4Tu3uQLwz8tJv7rARo+Y2ojR5zMb0fr+2rPlM2ga1iSXGbGUPvrxP1MRLlK4Osmp
HRrGfko3QfPOchPJZJUC31/IUtcbyLdUSrDSoWFMG2wV2r40UcV7HykiIJxESPSFDLGYJ6vN0wQ5
LOWcCX7O4u7qHjPzVPAJRWBw81E4dfU1a65xBV07BIBoFHxLAYX7yyKq/e0RRnEm866AJwjEZIzP
8MqAdLRjbfJ4hqAPq8Vv92mFNzkpXOlog7SKXi/hIaWO/qfEPQG/MCuS/FX8KL5n2XbgA0h3uJ+n
O8FDnM/v3MsF1Z/gLSiaYYWPxyYdo7Wo/7/0SHFDvXixG/J1pbwfvQkJPc2m7efb4V91tyc+Tctd
L8EAZ4cYTwCwO/YvO4D0ORVgSdakkOvug1/8NElpOHB2vx8/ebkxvMAWA3ZrqaP5YrmOcceeEHEu
gqs993EQigIn3U2KbWXVTmNn6/nY5idBWncn2kpDkyoqXaFNrtqT5onumc+xmlFxpjFjphl7Xjpq
NJSzBnEwOCK1L0t2ikcA0JXvi9D5GX/gne2IryfZAHpXh/AYnnYASFZLPQ+c/1gdFjrs+fU5+jtR
faxiOsr/s4aDWmrmLiAbaN4dj+Qj2/8awdTEMbpGX+JNFPaemZf01r5N91P0mIzgTPCRt5w5+urR
dPMVwpT7WX9M5QChAxBcXQZtEtrvoVuymsUYtVtpSlVmykEnWl4StiGLJo39O5MhsP9RNHmPvleM
mzjqHaBrcL5K5+Ydr0t6NRVPVlrJjNMpWaGG+TflFyfhKHw21MHPv0fLU3Tx8Otjq6p0p7JhZHiW
CTZmsKavJaEGCCOfdlBhiRPe0Avg58i2LbK/ygX0PXe2QB4dzwtV+utwmqZz7U6ik5jMmxmYKYkV
7cHWNwWUDTsk1uPNi3OkBRMSgUoDzhloFJuk341HJGzBOnjQrWWNJmqKVL5k2Z6Eg1PrMGtZXpuT
GVEKkq+hMNw+8vE1766K852CuaFbOUrDCw6y2YN0Mo84OlJoi96oU5x+/nfW2sd8eII17zwlf1Oq
H0jVg/XbJfNl4hoUWzCrl/7/GjvVuYAMBnlppJ7S8G3CM6tsJBJMfy1JNoXP6qR9EOzzXFTC8ZTB
5LQCJ3XCowHOJ9XFKWKLes/sLREnImQ3Fa3Xs76nyK0/qgxPne0zTxfjybJdeN/hN11gllvdedpP
op6eA6uhuUKDLTDoxqs3Lo5mELhCckyF9YjXcxaxxKNjHa38ChFRAP4mQt9lIt6DSXS8Qalbu1/+
azQ9qQbouijUq4FpAx22P7xZ5H/Dpp5s7UX7jS+Cm7lbPtEVWs6BDyP35o/eXP/0XUGL4oJwb6YG
8wTyn6+yfYcHrobOC5/J6VObTCGspmdUYy+yYX4UHd4R3vBkbslv1jg4qBKJ/sgTb3vgDCtYt/Vs
U/2DyN9VQXQN8udwkvpSarE1beuUXLHvHXBm+nMeo1M8vhPUi13/KrWRNxo3lFhiY9VgdJqONcqs
gTQsTlDktmHmXae0aZ2IQLZmaXEyEktP49bJlgP5fkVOv8k5AuyfKZVvDNPQPfgm/eg8cW2EAPXY
oTIgDzfmgedmaYlhPxAAn7NzaKCXNISxKeh1uj6bBUdR5551VpYQmlHl3jEemv+A4KZWQS6X4FfZ
kyH23eaR/eLWdXyK+7TfydRez3cteN6iqd0YFj5qd+LyYEpafiN6Xu3HKfRIA5kuvXZfKRnSTX2J
egkoIV7grmP824mF6SZUwGIZVBY+tIyRdYpa78zcdG9l44FDFME6onv1BihPLehekfSOkE3hYbhE
o8uchGdn/tRykGH6IgmhAJRD8UV+UCPYIV3iTMuguGDv+YCcYDUiNkHQgRRqu87wkq/lr5muxBMm
4XRMdTyiKxzlfsG9o5fipEVSUHKvFWMC8IZRfxZ8rsu5rZ4ywbSSeYDMrAlbBeMtmx4/WGlyIc+h
lQfU/+zVCPI6Oz8fb2/vdGc25KG8ojzOXOeJDosMb52u9gbHaF9HwTjTAemnWVkd5/pb91kqfShL
oYh5Vq9Fz91386af9tv/TibJgQasERSeLDYHqqHp9zBHNTVEArBaIhVZ6R522GcSxdzvN/IxFYaD
uteflaInAsjRJA5q2ZmbB/s/UHZ8ID4whxMRyd1Vk7FIbOu2IAj70jTTllI7TtZ+YFRBADpZ3Vqn
OkFN53X+Fwslf959BMFnyyZ4udmhRSzHUMiecJwrpbm3KG+qo4f2GZuhTG6zwl1m/jspDHHsoISb
ozazZuJl8gd2PWksmUx2Iq7bIEnd7KvjsBKjTqyQsViXadahUO0UFIne3qkXDfRxYDHMLVsvXLLg
uIJWAf9gS8UZtyd2Ef0o6LwlG45dTAbM9ccT9Vas35POx7IDrgvUXuAb3Lg8H7hgHPbuxi9cJ7vg
6JjaSGH545UJSibUrbdN0WBPrR6gxTPz/nWF0D4tR6wnBtYIdmV0Sq+Xvyy4p8l4taYru67diQIT
wvXxfW1cEkhF1Fin/zMPV3YrAwoAKMmc/btGHQyC4DlpZjyX1jRdv0lLpOdgofAhJG2JmEQBifcq
LECJPH2CmLeQH2v+NiT5mT/gSv44l5Jqu6cyFPS59yjjcsgUgDFzCRM6zCGUBFTvCdoVB8bf17HA
t3rVN7pLUBZqPjNbi98dfVOTaYq6Cde7E+tQNMhI3923k+6JzXpCkhMRCw1Mzjh+rOD6O+RyyGy1
Y2BUF1T0O760TkDIOW29fAcSwCGxhluSSKEb3R3Y5yZ9zRpj6ObzCQ+B5eVSTRpGMWw5C2x4dGy0
wyQKse2hnSoz2v3mNyOdRDwzXKpI96gahwx8j3iR5DETBSObVccKbgBxynRRoXu4Sl0hYJYX6knI
q2e5V7omQEIpICUU6dh1+Jg3jXXfDHf+0f0y/Qk3qhYe59gOxamSwBkrQNTGU85WMcw3KSRwwfqw
BwEiPiqbydI/sKyjfiJ7nv6XOCwdr2JS3P75gFhOX2nykgSNoJMfXNBKWzKLklIxGR0AHF9KLFvA
jCNF2M02BkENcy7E7Ojtvri+aVorgxUeQ68H4FsWAs8eaXTaSrqBqrP7e0Q4MOO9VXPpIlSKybZF
Bn1qVemZalku+vAwXNN1pJE4wWUh+3a3OZPR48Xf1dF8KrB4aNa7Ol5/wLjr8ihX95dakBozsqLI
0uXGgHGoE/KcqYTD+HIk3pVGpUylKQm1pRGb8B6DAa+rdoGQ1BkhP/guJG5f35//yfPb0gWdbYNz
ocQHHsmsUeNNMSgT9yWg7m1lf+JmzW7hLaZ47tliJ+7ScHNZ6KSjF6RIgHpM5H3Mpues9v92Fcla
7CLX6fyJBMAtHCb3uYTX4lIT5Vdoqg0MRGK3QSwQXOHHVNkesJ+jSpCZupA6hszQa7RqA/KE8BQm
F21m6N4aSVQd7wE32QWlnRtnxL45y1sMvKKQN0aqMKOK0k2M3QwCeLFysD/XZOkYkcFuL1XyFpty
0FmtCgnEQXHtgyg3tiQ0p4vnkVK6ssMMpsbhtN0w0wYiDHEU1DY5QOX4m0bY/GQEG6QTZA8+elO+
vshuJA8KHOAyWaUDgKI8PD/OzehwbhpBiB1VypuZUqS7X7hqfeFSkeTyMm5Zxz6v0zvXHyZ3meiy
h7RHqez17QkXJrT89IhDfYZfjmL0c1xWNpLee6H2J6e9xx2i1OiILxq3neBS59PL7jAtKFHykl2w
Aac3Yhmd01vKEyG+Xy1FaOuyJZc0XH1donVRMsSYutRQnsfhP0CrIRehB66B8S79Fur5noM/t8/6
V4vuRfuPOZXCuhevEGnowL1cF8/DMeABTao0fw2ljNNow5pgMYDlZOmuTrsek6AzssVKSOA0vNhA
Zwik2qMu0RWVF8LOO2TQZzZW5QCFyBJKhvzDtT2J4kOoSZ1BWDKilGOne9eyahDI5nINbo1ucCgk
k7WLzNwMPe0HOGkmIIEoqvxkxVO8pz0X+UUyF2fiOw4lMW26gi7rApoOwx/R85TkyXbWmS6ijnT7
H9dyuviSaOQaz5FI3ZhUMqtRe1Or5tWsWedPfgJbJqwfHkmebM3samgc5qLkls+Yp1pTYbfzaJ6p
0+m9kXsuxwu5yumrdVAF5mxggIEK8vD4pL8pHMPotQx5ut5DHT+ecnSUh+EoD1cY4hFjGqGqUzQT
MQ821eKS55Vyvo/ChM+gPavVDdrg2rSoBygQ1VrwUYWWlY7/iNQzgTiMGYZLwuPZBz/xaStA4384
Jv+Rn4dB1KmbjSS4YjqZFjATd+w/gtME6qKK0yEbNPmLczwjN/1VjD6m1JNKvmawrblKtYyCrWgw
hgmj+QwkvavjCxwVJfmQxPgSF5+cq8kVvIa61EbmT5wrjiNReylYWd4chBalldAMowjFdGIt+Z9A
45lJ5itf2Rojvz1+FwuEzI7hrhO40jQN1D4ea2LiFmIFYdTYV+DcLDYi/Ud3cXHj8RMJar/pZ55R
2g4mGpaGvZWiLEfqy6lQUhLPXgdGOpBgYKYyZ4pVP4T3XnE0aCZESz/8YZqSsZiSOWO8pwWbSyJN
OGH95ZPVNXAIxL3Hv1Ti4rUnwyrm92whL0ABHoeF3/8326gjw/F6t/5V/4gKrBeWGQUicYHf1PB1
LIN1rDBkFWxmVwMPm2ZVfPPLSoTuDNh5oKDbzUq/aIQYJ9OVXo/QfTFQQ14vXZScWxaqq0ipWMxR
coTjLu2aCyiSKavlhuHxielpNfF4DWIfoYZ0NI86AqO9vmZgjN4gTpVEp45bf3kDXyDRVb+lnbUd
YCQ/TyjHtKdzbR8v3MZwC/M4vGKczFa3jyGQdgoOpdifHLfpVnNDIiK0gJ3JzFI2J5ZH3yXDh0IO
ELdKauwWcpBiqABJge/HtRM5HYwt5PE62ecw5zlG+i/mJHGVDz0w591EfBJPqaHTRY+WAkXdCKif
Gv0X2chCLYAUgeItq0V7SU9BRkDO4jNw/RI6aXeBoaIXksfdeNIeA4yQsZVNF6bt5h7B3ebupXfB
w6vFG+xsWGQVzWdZSZ/Bizfoh1wltwGFtzSV19lVJ7V8plN43KkRLfqk40JYLRBsU856D111oUi0
ldnK3TxT/LuG2Ps9x/lB0EtV/MlOw64mv8wRaPZGc3Gb4yD7T9BJmKb09npq5c7fspe+u48fudDT
7eivcb/NtFCXTAhT1ks6ms+bxfKLLofPxaVYNS7qGJsbqtXB9euqWlGEf1O01sPzoy7guNv+hva9
A5FC9+JyjSCdYQ5rympcXNICymwEqo9zLlr16eaAWWIcjsITY8yCvgQeiTQNYml1hTmAu8RXEsEn
pbLrFiqB+gxKEo7KP5eIZTT2QKSQeLbpdvnrOz7mvFUSW3xbSqqWjUDFxrZ5TDWMHUC2WAZZ27pI
WXkCLq5oJMFfpdLPzonHKnIIw73gRmGuDFFdQZDiOE3UHEWDL7KJSq4rXCZ5KA/1cUWDXlc8Yhq5
BX70AHruNz6HUASXFDJ2ISxYJasoWL8VICDU3mhl35qCl8EoLpIKruQonNIalteg7cq8XkMyIqBf
Zi676Hg6FGjKYS5VJKRymbEVJE6MQ7dbkFLaOG0Luu7nIr+DXvb9YCXkd1bcCrPz3cJWoYw/A4ed
mV0o1jxpAk3uw4jtzfyozLHyl3GtZ+yNSAar+q4rR3xnPAwJPazNmtOeUmlpDcG7v6rtnZhcqY3Y
pUTzAhBB3pMl+MdX5/XXhu2AIXHNsmQRZKC70lLwd9ukI38ZbOtd65cSWf6oow9hMHAwCaytvhFz
Fzr6wOZNAF0zJgoN+c7v2BIEqRwal794FLDOLz9ppKNFLP5q1Ohj5lR0MwA31bE5QGKbtH7N+7Yf
JN+z6fArP9+D+picHXVpHGDQFs4lbJ0JT3YV6QWcBT3U6xFV0kto5JkAy/pD5Euk4fHukrPfVfrG
7B7OCaiRGBB2p1qYVzx4yeIIaAZcj+gh5aGjZLcV0pR01hmXE62nfxJeDw/RAo9woXNnm2m7Keqn
5B0Br8X9hsU0MN1irfMNR3pc12+PzKbqoag/gnsH5IDuBTCW6dbamZIyZFT6GWDeDEjDTfXDulF7
HLpREW7Z8NVxXuxIDbK3cBi3qGBaEYGMRsOop5bRZzmrGDYfZ7Zmj+tGVDi2e9+iy68VPODJgu+7
RdKtg02PTB9wc3iX4dFYaWr+9j/+Rwvi5rrU9KCzPXBNEkbHxFNPGmVMJZjODFo2nc99MRzODfvX
Zqo8EzmFP92XVryyqIa+J+IA5UJaZdKvxtLvygTRnc9Dex2wG9BAjZOVe4R8vWhPWo8XEJS4vyPo
Z7EapB8YCfQ/+dL/uOw6MG2s/swBuiS52xG/kPBNYCyaOKrd/reKdJtVUEG5VDzN+5rF0U5Erfoq
ZJ69Qd/V4HoUP0bQV2PA4aKlpKOLWCeIodQjfM3qsNAqNy1M+/Cw7ZAVYMQbpL8CdZyluDu7dxzX
71nDSpaWZGW7Vuh2Y94RsycKPugMa6nyVFf+PozuxXThTC3JWqYbVO3lYmDGROEexeR8PdOMt5m/
z3KifPEyIeafpD+LmJqRVShxpOIeZ9LrB6c5Alo9bHYkVcZwsBwTvJgcnwHhqtHVSV2/9dxSAAzp
vONP5cV3ZcyASVP++u/jmWoQOjSdmBrsq+blORVc7yxHiaCKIVPlLNywLzvbZDM4tJyJfPwtQC5Q
QyrFFlfaKRVAHfIZJ2iZ6YC3bVvCd34Lkb7AEQ3l/dzzQUEEXs/WC5zghjPNhtro9zLvUEyjsd6L
h0H09RqYmvN+nbyNR+bi1BfANJew39oVu1Lb0ycbVLsvCekCV1IsFXWIyJBbys9MapnqqVgQfa6z
xEE7JonVe7OkRKBTOY41EdtWFaPtF9G/YiCxKjl/Ai0pNeA85H9ljr+VQ0SrIvfwAM+koajqeblP
+o7lIgtPQ+m/7nKXDzVMKewo13VhJgwKY1/M/Wh1Jhs4dzDTyl5AU+Se94x0AL6dtHwrUncTjBNM
EOchxB8+ZlKQERsiGkk0N2es5LeblkxGdAem+8UCoQchbDxunNLzson19eOLDhbilzQOwAW8O/BV
f4fxTtW6ttfsK7osooMxREEvu9k1xKGPQ/zDRF0Mf/69yKy/s7ycVNIcEHhT3J8HHYDrcE65cLT2
KuivGr6YoVzE4s2wRtFxMCcEk7ISsksUYg9uIqNM+DWOOqjniu39KnxxHNsjnNB1mPJ4GFmi42Ti
xSYOe/J3mqo2fS2cBWp4Shavj8aingoDstOSdFWzgYcJgACitY8vcAtMZjiqg+O8J1DirdmAcn4R
ui93YJaaoTWvN7UIyXf/9TjovO5fPTu8ciZ1Qn9iYf68XUnqtjm5dl8l3NAvQBdq3eJv8SivzJ1I
OpCeam2tqFw/jLInz5djGk2tIyre9oKIo3yLod8sMY3wXCz+dHNHGHYBiz8qEZeIyB3f+EcgxrSX
qkddYjJeM8Ztj1+tRktaVLmXFIAB4iz8MX37P6IIsnumzu6DU84n/tWYpa+98wjoqvpXldEy3XXa
OgGwnY/THaxDUicnnghmgTQ+/HsfOjRdT5VgrgDg/5o+sX3/1w8Bp3UavBRNj2ojzQHL9cZMYBbT
3QiDH8EM/ov18ZjnpdUkjn19MwlOudsdkke9UA6HuvDPz766lJEM6KbTrMJ/EpFRXruiGfm5bcYE
8Dqnj6pdIIbBBkR+V1304D2ciB8JvG7IUh+Tv+gqBGPvY46MdZr+UBW0PrAR9jwu6x4hO8bFkATn
NfcQr5YCAXCPuQT40ctjolK78KfcuIjzoh2X4eBpc6Ju35+tkbiKzq7BSOx+sBo80tRn26nsv5ck
CkTmbXMBDI5YhuEJvNlSAKl+8sIT3PcdC9hBW+akkTbyStlYCC1ocfFWIY8pdpDB2sO003EnDANC
dteUYepmXFpiAI3mVz+ylO4QC2+ElPQeRNNj/ZXJNPX/Ce3pLsFBRxmUXBYJBgEHIn+QLAS2s/2y
5v5kbo4HaLYRNFHIgNCT5nNWLk9UOd/jFWivq1cMkO0rnM4XjZWCNuvRDv1Xke875XakyQVljqsr
5vAypNcgHTqoLjX7Rcy+tVpVsDrIimwOKAt22GNEbcfwvaIcw74v96mSeuD4mc/j+A1FpxT6flg7
8bP4j96ViahLotedUt+iInVZXR5Ya+zEHGKJIcMxLzMiENKavsJ+4mNTHCo5cG2wOY7fKz8aMqMu
/9cfjD/fAWm8ggYfTzghzL6fPcFJEDQ/I8NQQfBbWZcEfD9okEXtRIJG0MH7FAi2B16EWoa2XSu4
RZ3lm19NyFQnAd2xXb75yGT/cva8HuCEDWOaL67acGrarHSOYny13g/wtiOmqjXxiOLg3tzQwcY9
08QU9/S06Vmsm4ykfb+Kscn3fSsIjt1Sz9kdzL55tIRhMroqRITesj7Qe8sGuQKIQfBZ7BR/uREd
2wDKi016Q7LbGAmR5lG96c+VbJx0cI+lZ/kTm7au50Q6Kl4bxapv5k8KPKwmcrGcDlj9+Sk4Ttfi
0GiAobbqHTtazSJ/Lgt97fokJtgpPZycfqXcRjcgJlWVIbMQSUG0L7wsOZY0Y/JVOmSxNfGt3Wl2
4W4GP4znZBLKSZWn+NgWKdjSnL53qhgbLvwYyNylw0z3oYJCRnmxEPKSg201weBq9pDsISCKoMOp
wGm1VnqPBnqcFsCsuXoIM1e9C5eeABY/TSybQvg8rUcbbsG9hozThwUzAw9PpaxrxKjIBUNu5lyO
JlRKOEOYoaJq1dAuUySlBFuT6aIMbmbUGvKwIr9kceE5EHgVQ7ItqPUPhaDNE7I3b/HNrXfOxVyL
dqH3EBWqMQGeUqlMBRystfpP87BM7rxA6Of/ZurICOIDb/c55qei/i35u0XbwxSKtGXR1crpFX9T
YwRCcjCgI5yflYNAYVvshgiPrhRM7xdBvXznzL2bjx8j7vPEAOoIonjY0q1+TjkTFB7gIoEA1TuT
VBYrRhyZrd8Kfsg0/JoYJ0nJ8O++km1IvuoKkjnQHFurZJMrJahvT4ea4liSiR/W7oDVcegSqKPu
47ff0PO82ARWXOQsf4T8FxQUFKZy4K+D9fHmkf25VRsOmlzQMbWqMvXK0HQPjHy/M3zeAoF6Typk
9O2GoourM2IcbZG91BfPLSQ3qy46tWqk/5XlldcsywC3OtqOLxP0e27NUYS44spKuZ/dPhQHrPYR
TgJM8VgY/mu2Rx7nWvhPLfIdOSOd6V6LYYSdKxKIINQnobAN7XN3dDE6urpdediKL/Owwxq4qMeD
PZZYsGzrrskE++LwHQJ+0qTy+coobBFPxgh3HzpX62ti7HhicrVDuQhuwHsu4wP2SVFJoTZUggAs
3eF88B2D0eXOL5/pUgsSoGTqkYuH8sjuLCcrogGr13lS8lmGVwxjqDOI6Bmk47PsXaJ5cdSsBOFN
0es693v2YD4qZUwsdDUmTbojEdWEl1q569H8ZyoocfDmG/WrObZNIk/RXMadUYJMUhZaJTjwwYhP
FUFHBnFvoHtVPQJLQKmW11skz2zYxwNtFVkg9Pr5BNrldDyGN9u423Byk1C/w5Kah8i7bBMmAMtE
lvtFzTCp1SirEErQQtzt4f358bzwM96LHRLeV3XQsyDJ+l5lxGZz82etrVegslL62VXUFHs8y9A+
OyLVV9ptFzHVMlHd+QnxCeZLHajI3Ft/Hg6NZtBGlK/xtjTFaZBjfaLJbt+7Iu/4uGFYQc+GsZUQ
HM1uYv8A34W+0DXZAeSjlIKwZKQZUg00q6xYMlyWq/VLHQDTPRi2ZPdrLepsJxe9zT6FWd6iFbfI
uwsQLCz8tYzgCRCh+IIdYlOzPbTB/GcCPwO6w5U5mlti2x9n6RfEzm4ygHDHm4099wfdS7gixav2
89Bg4r9iaHhQHZ08PivRnP1BaU7BZuoshf4xe67EU5Kfsl5Tyw3ZmnoeQq1m/iQFGUz/YiHyTJYm
zYl0NrgLyWMwdwUqsdc+WTYyFOQ69rahcQDDDIb9vy8mvgIy0uo9BWZ3kYsx0Y22+KN1SRDxISfV
agXkVvxOYmcq5F2RUFL6KHnKtkl0TXvc98OMaJer2a2PT7lkYnKjvoKHQVh65mFGHdO2422nnPTb
v8zh1Y+60gjxM9gGfxQL49cnhfnp14vb9Ag4aSBQgzUABhHh4toufh0fzmhymiHNismKKo3GYGMc
sVgvad9HPTjb0PBirDnm7kx7EDA3OjTT4g4T3ESMio3H3or/YSqTMvABbWWOEf12EhtvpDC+7naO
JcOE0ltrcq9Habkq70OPZ3woBwwr5FM3jFepsNrMEsaZ0bcaX/V1RibKBi+xUgb4NGCT1ph5/r1V
evnxdNSctGP+hg7yipxjNkG85E2BFKtI76cbgrksnprXc2OtoesSbfqbCfrc62fu/mVXqY9bd8tJ
jNerUWaQd5bs1h7xRXZx4+3qh7wbYpeVt4kWsWq8piX2sz6kUV6A8aRetyUdopH9v1ktk4f8T0Tf
06loJJeCMI8Y/7cNL13F37Vpl0xHaYFXWDmiC13AiPNylE/eIBxzZL8A7zflHrcD9XxUgG9/uVzA
dReDvvDGkcyrxZzw/koobhyy5cWD4AZD7pfST30d6VDkQAM4Gbp9K4dyQBMRLRIJDUIcMWLJNggS
NWRJFiz5u/1mLR3wJSrzvAH5caP8p8dnFqNBhnFKKrAaT4ZaIekM20Yk4LwMHWKsydfmY4pQwDpU
BVXVEaELFdIGIJSpWO5PywfaMN21Sq1cDSZUJMNlzbY0Jth1+IX5YKLKXBUjsim4BhPE7vaI4a0a
dE7h7zoDA8GPFmGNw6z/jajqsERk7H1ev3wNLY6FQJGFuEjmUUUhQkN9XMCnISbAkwdfXF/MtIeo
9Tz6UDRd1V3Iyx+k0nD2nJzkwy+7NfjzZyUFwC6cEOwOj1/6Q8X7KPiO+CW7mhaBqyZI3NDTxRld
g1os6/cNAsrWp8WbByxuan+/zpAogOMxELw7/ztWNYho1fH1G/JgJ3CQdU5xthj5Y5Ani0d4pyeK
OzPMuhqHJoAWkHoeT3qHsy+f81FGtB+lA2/xOu2tyUUahIxXXkKYG9f+uSMNvRccU6wYu6HnVHdN
APAFYz0mn/JsAwCiDHuJofx3BiO8aiB3yRWGsCAYf0MxyG3cQuZqKespl23zsDRyllmCXO7dA9Cn
OFEnpNpEDtCzw+N8pTj3YvHuU9azIh/YTqzS51R74qn54gIUE/W0MzWOwVFJvOZlMJGs7F5WRJ1S
m9iTJCKaSqi2g/Hv5B2scSVaY4Kiz9GrSGKcTwQxEoPQ1FnBs/oCRqRYKj0dLcwrDTVRLAax8+kD
jxHqhdeEL2FU1+xc7N4k9C5ePqymsaSRVHzUQK0bgr/SbpgCR6dD577h8PXu5RiH2KMQf1aPr5sP
QfejKw+9fculht+ucJ959vkwgJXNoAW33cn20CCYxMhDKEq8Uj5eA4KYZaKCUR3gA0a3GaLejuNx
Q8ogvgCbjidQcMBwAm0KJDMErlT5zdfeNHGYCoayaCEF5fWZEGstn/S4B9Y/xtIboXGD+Tbafcs6
wN1eNUzFPzhJV5ZdwtrzJ1lUEU2F7jxUL05XgZKV68SavclVa0r0xSMDifBTTnveASqg/fyDq+JX
kevPv6vJ4UgJyZLUTPrUZfPpS/cAQ1wKu4PX/Wo/nAvNiPdVthJIikT+Ba1Wi+RIFFiHM61hMMcy
QOEqPRE9/31zIgweaWztQRo+CLifgBHt2vgjyLwuF37p8F4JzvoLNQhEnRdeNLrKRUraDgymGCF1
HXHRt+vva5XOaR5Q0FbANZ93zPuplhrZa9b1WUfsVxZt8YnpykjjIW7loKbfRUyYrgoQ0MLiwud0
o4p9aeGVgGyAODFnHbkWs6MGsHAxDe3rIPjPAVNsD9AZ+hfq3aEV37+LJeEtqZAPutmUIuafM9q+
s2dNWO2D63ckkWwHua2Cygz8MyqabrJBWyDbzsm3AbAjkW9NSY5Xg4mHN0uzjsaygR2euaDZYnKk
aoKeMxVPEphDM5Pc09nzVX9Jvljsv7QSwhQXmfWWcmUlGrPCT7gGt3H0gkqtNqLxp6KIoLyvBoJ8
8tJWeX/1fEjQmsd+9dDueyklZ1SsZB1JI+7x+3MPR4ldosSv/oLsPE/1EmdeLrAEzg7jc+ejL/bG
nxpEHGteixrR/TOMQ5zsQBr+y3kv+xm9K4CLvANfADYbyyi7feQryWzrVn++rh/ybtsCO1rYmUVn
USMXUPXsmotmVfLSC64wrkp4ipQJJvkBy/1zAcbyYL8FNaNTIkIWmBz8u9HE0yuVTq/7itdQH6zB
3JJYXwMJioMI3I4FDvVNKfd9YWFZeWrFdM/akq7VwOzYx334BiXWswcckavcIr0WNWYKfENFkQVL
KDbE8o7Xtb9SDxL8+/wnRWXDtDlKFa99aOkRxkMPqSQqC9vI9wFG3g5Ktp/q+aw80Rqkb/38E9nC
9kH+q88iDgp1kJZO3tGZWTFR7K37/ySJ0tesYP5ciPvkVdRwj9bSR1HS03meQG7qaExQEOC1tOlJ
B9rc07CyUlMsrRXFhtS4d3LPTvxYA8GubF1LkwYI/nSIyfGV9qXCwSCIn7+3Qi/1GBrYFCDqrzlR
yRikBevDaCy/DOk2WqDR5s+QWzvfAuC5XTScLO4ISgQKMi9++LoXiVe4e1KaynR9Pd7lZBwD+QP3
agU3jlTXlQr2DPfpa0Tk5dJ2FL0hnlyL88Ll+Ox05jrcZ0wkYqKniR55s2o4j1Ag/FDR6LWAc6Pv
PVhkbh3S8DnuADqnJ9geVK4DHp2qddOhG7jCNqH6Yd7W3NhOGzPqQIEqyM8h78qTwMR1/jWbIUDA
Kbhzs1zIoSgDyFAW4n+xVeTGz40QdpyulePNiQxYYeBgXbEBDgDAGx3hYLtNlRJ0ZbNcRFgpbCLW
ca3g17RRhuEaRVqcBXGo54waPQY1bK5yC/NvEyAdK0K6YPdFmYlZK+sRGMTYPNvoQNB//J+W5n1i
rERO6FDsUaIgFRz+WgvHfFELWLC5iKG9DW/uO4lhLjGLafdoRE5duZxZZ1lWnJo3LQdc/0VMgmS5
3Wu1OJ0fwT+xpwb4fwwojbAqS5sElPE/dWJ3mYK7Avbj003IIsJxUJsA72Dmb5WHUuoeCtbhvGAV
1OvEq4lS8G1vqje3JcAMaQHhe0OqRE0cWmDREmUvQ0ooAekHblRF3GrdH98r4qR9CCG7fT6E7FCn
povpJCFcX1GagE30Qy9fAEdcpACTMgh2n9EMrnCnDHIwoBkF6h+4EBYQ9ldSlwj3zT2mDyPT2kNK
rvz5Q5pisZgQsXttI/FGmQSGPpGppk2nJaGRyWJFcLa1nh3f8/r24I1P9QdIeHcXGvjXfyKi8qmg
1Oa4dsSilx3S7eSqDa/QEcpe/gRt+kAd3/BCsk+ODKPBZ6Y3T7DXAXFoYHQxsXXMmkma1Fak3Us3
TR1rGg7IsuC39qNfuBJmDfaottJCJeoq2NMSsKpCZdGBSySq5TOu6iOz8OLbvxLzEsTLEOkdKZTl
wWEi8CUm/d/mLrV57/+KoKifgsQOcob1Tqgjxi/jk3s58AXS2N5Mqr3ItCubdVlItV1JzsVGqtPW
cXf6AbY4pFMsdy40jn3bAoMHGie+Q7BZ+bt4rz6E5HMKIyJFAjsVD4QDLm+/UUT4PQ4ZPlzcLxD8
cOqHkMb8k9WrhdRum/V/Tb9cCo+t6SLXsJ9yNEqBvmCyptN6XUbm1aHwlq3h46a4EMzT08HyK08c
CYKL355FPupQkFWw4iO3L1r8kFRXZeKQMB1zjPtT9mMY/l7NID9iCc+GK5kHku/0w565IqSOP9pL
EKEEGRq8tqcoeEuc4OmIAli9PkjtjUJbLlH1nG/CVAy9RvFZ4jGlFBn6sq+p9pMyzzzN/WeSBE2f
JcSBEKjfVWj2kjt+Zjjm80nHSzwqXp7uTwl0X6ugaFAlnwPz/iJfsJ98dxKfd4zLrP0ZddnCYBU6
6WPxRo0zqQtCOOdmLih4Ux4cBGzPVIDgdG9253X5E1gay8Ho8SmWsnAV8D2oH2c6bROtr0P4iidt
aWJGIXexjoPM5Pb2UfNXOUlaj9chClSckE9GMgB8q0KEYeTRiT2OoqKRauXfhm87+VsKrEuqQAH/
qsYK+O1hTjQmmZ9V/EtGt573vBNYIyJ4X/qlLGrPqUJE/PTArvHRQjKOk+FLhf++5Isd+DwMxOmv
nvnIlh5WgsXicoFilP7yNhrhTpzcz2Lyn2oxE3Xx1Rz1H7dEt3b+QOYC5hcbOEO5YuBJygohcDdw
wPhLgOBviBYa/52o2oJWC5GxN43ZROpRKRKc5GLGp48F8U4jOGmSjTm+IcpH0xAHRRn/FG+Y6PjA
k1WNMwrvTYbTCEYVv+Zfq9ayOlI474wGD+zfpixnPnoYSz58rLpfFG3zYUN9oteSJikG3LXOoxyJ
T7xggb/JAzgzYQSa/2XMCPRo38US7H7Hz/WFiwiK+F4pPt7fXHd5mGfgo6Qo7MWnct3XMgFCXcaU
ZiiWsa/uDwssctuYpAS49e+oT4Yo7andpebNr+2Wxsrl8ElrPMQUA7MGQC6MO34FL3l3JhIgA+yY
v9gWd5eodS/Oz/Fr/GmCtJdvEM1beSHJbm4uKDvCog0+PDAy9vfPF2Oss+9xtvZVGXcbJk78zu/F
dZFepXfHTJRwSCjO5GlTZpd0mo2zXsw04BG7URTjPLUJKt5sukIUINL+isQXaIoXfjWIv2F2rr8t
faViPqWyWx4eCjEFAjy8ftIL03xgxcAvIMPinSxW37VfolXoKoUiGmq6ppNPxM+t2p3o3OifP7hv
V1P3NqGncVUdaxz6891MgrGXzZ370V0vKk9XJwWd5ZUFZG24oqB5qtco0gbfGiQSVy0/3C8Vvuvj
vub4tOGSdko8o0oPN9rCTRpC+1r+Kk0U7DteLblxn+YIMIvL1RbM1uYGVaT01ZmHVO2DkVR2ULNW
bKIgMdD4Dl0Kf8YPDdwLRuyMVW7+Zm9JL410oEFGgmuGvxIXBWhDxmZQX7bCfGteewk9FF0mIshm
mmI85XXG6c/vzLaJ9gE/Mmu0Pf8IrgCL099tUPjCBPqE1t7+kldiAHpEvAnVHf5oEVu3Hh2oH3wT
a0TXM13RTkKr7wCcYxu1hIf/SKEPNyxYwJxbegOH3TWOPZzpp1ZI5Unn4HDQ9+0MD4t9UljB5Mgx
0+Ru0zCgqNuYcmjaONnDxTGrD/HtvrnxQgIegeKGU2PZ4FC+ayUpZ9zPRVieLuLTdVjJa2NaZ5SS
3W19SiRLN+5FqDoaORLdMBB2VBPTgLZMjfv9WKCkveepI+m1fqfJlwTop/IjW5KsLxWdZxBYjQxR
hQM3lgcqkTDDEKRBXN3HV/vz7FqlhpZhEjzmJF2I8s99q98YuhtpC2Gdtinx2PHm2Sj0/TrdmCQi
yHvBcXMu6FVhprrO0K2upEraYoUxkp/ycPZvfcaQelYQbYQCrBQYxcQz5iHbx/0Ozx7kjlcF5gSA
J1g6W1yiGspLPBrgkBwGtSccy6hFpNVI0/ggZgEPo3d9gdR6VzxhyRNqMgFfwVftzdgzttKRXXlq
PLuG0ztOuWJ6E8TyrPPwrWTORcm/dW4LPDtTu+xwkLG8z21AQmjOtSvI4qSqqYXkNYPU8Nw4GKK3
6xpvEAJgnomXve2PQxy+4h4GzZYGxXiQ2jyWWYiF4IjVnNSq7hXgwKqOxyNGlO4kZn8bb9MX0aFL
+rBxxJoHTZdsdYdH1Ef285NjXGGV3uVx3h56N9lMyMeaQA8SPoSPWSUJaGD8h54oNdbPE3l4cHH0
VzhCnRbv+FYFfbpkVFJZtyR2nTFpe/ijDbD5hmWrVcK+GATYGsodWXDRjQB2Ffri8hd9w2iGWOeb
aX13yUvreFTijY4x+mSJGbVAJzfA9tP++h1ysdr3qDCaYz0zbtOisMSQ9rilJ98VZJC0hzd/21H4
FZhyNUoxNsboye5fi1QekX0GKo+NIc/VjfZux0XmBVo8NFusBRdM3OYCTzNc6Jqs73lHkm7VJnLm
Tnyd49zZIs2HY2DmuO3OBmFvafoa+sX49IuFGPM+zecFsZ0P3yRb2mSrO1KMtq3XkNLv94jMRsTw
WNLZUwaUmy2cKtqoMHi1V1oAUxA63TBn77pCcVYJPTCphvEpEn4qCaofeZrJBebtwTSSbfseeE1o
FSbbcZjzGhz2TtEiHV1RrlMIxuy+6a2S3S32QUVz//Rl0gAp/XKCVtom89akBH1ytaseYd9bGAYV
63OCBC+/9zOqC6/iUoDf40bnTds2yC/2VpyUizajNau60i2U0+MC8HHunxo/trqqdkW8w0VbfTh2
Mgt6bIhMbmlADgKPj/bfq1mbH+ris0yJaWiQachej6xOyZAk/v8OjGupguekZElnZ+eNezYIFXOD
JdNrz1Itd15vp03MgBibx4k5IuzuQFqcfHVxZwxT7Eavy2KknHmMAbKB+l12hTGaQ/rSHprKFe9t
P4xXeV9u8Ipo2UZ6VL453cmWXqztPJEKI8FwkAzV0OfVhEMqXd/FgVCSeCmX5+7cmi2Z/UR2wzjs
KcriZtA1xk4dycZS47bMmZbplwpMJh0Q/aJs0dN9BPWZkX/JGOr4CgQlsCH2Q+ErkmimsJ9Hxh+Q
Msu4ajzJEPiPNBMIjndKL63Um3j7AXYAbnEaW07a62qC5G6ubLKNWQuNzX/zrk4Gks7qNQiiN+N3
REiLHtaXhaCY6aA1F+8527iUoQZDT5DXTpfcOWUi1RE+TrzVA+DqqJTJEUrF0Drsd2ve5GFD2fup
ZPfDY8DuHmgJA2cQpgsVFVV8zesWbxuRkRxQmy5R8IbyFV3mxrrPrleQD+Mng+H3BBzglXZBbe4J
G0HdPM9ztHQ1VgaQeKDVE6yTd7gtzPzBMX6CkIDtjLbKElJmvB4/vTVLoE0L39tC652UIolTYqsK
DSWIWu1oweXQkyKheCoGSZ/Ygoyto8le9eEeDzZFFG53xdjj1WhnoN38f0t6LPnFxBbv4JVYBe4+
/TiZ74eKaQLKn+TK1+ufpvZdVmW7xpr4i4vTSc0VAZl/CLw0+C9g+XR9xKSfaHBsKBQrHzwzFuF3
nw+cxm6pBDJjFKbWupiE4y5EYMg/gm1clqYIceYnMyiAt12tnWK5slg64JDAD3XsDbAvv14AMGPt
2Mu1Qnyuo5dMjzbXs+6d8K8SjgkhzLONxShUxjfhBVCiZJET6g9bWQplPCp6Ao5VTGFQxr50VqNN
ah7GoAYk1RPehC5lZqEEr1wsY0lOCRHWXSqmbqs8jHFgK22XKqCQ+pF9vO2GjBZnQceOyKHp5eKl
ine+yp8sVFIPBTZeJG2w2osy5bForTPf8iWM7zgfu4evjqWZoyBfFdo4qYDYvsjsTf1xoXtFUcn/
krN9MbPZRBGDUh7WPKukOsD6g02M7oS5bEIYplxXsbCWxKgwYT4Zvvpjvp0gaI3Of+DKeSJEuFJ2
Ffpu6NKCdNHW8vHM16P+NwDKh/UQxwr5tOlbFG3OwqDBK98B5/EBFGPZGjXqhOC3sgKK6KTJuOda
us6WUpCbHC2ljtUxD4Nv6PdQCInJmNUufjRFzcVppW40h8Yj24gAP7a094je0pJ8xpLiKlFB6HJ7
NmH4m7WjThv+szrXIX3H6a3ahlx1dyw5WgdmQIPM5X0chYB83Y9aLoglR6W2IKis8I/tloFVKzrh
EqDmO6WblLSvvm3nfC0jqLdKn4u7eqOhCz3iAFq+wV5hRfkFmuNuKeRDtsiqwmV0UDAwBwBpQFwe
sF5ZVO8Qtnqse1NXFLyTh7iKTTrLlsJG+cVic8xpI3UwHoHwjwaLR7qI3qRG24CLLm2GKEq3C6QD
vedQaT8gMQO234Ak8YnVESikZSNSAxDeXn31iJ3y9ZIVNvkUpbG945mFySrF5Fqmb3jp9r0arwg1
eP2j5q2yyU6bsF43MefApScNeQRd1Hv+I5mFbgxddFpYBrGVleW0VYtjYTZYDLPTNGNF2vfQTP01
dP7yNeJTGCDtB5h1Z9sUpm+I3AOvloQM6jHw9GNxfeRpRr6ZvD0kymrAjKn8+IZB2hA+6Tzzq/0N
T6G6THQzoDDHvdmzHBfaWtO/m8lsUqxj8S1DtuISeMMrdx3EJ4ew2Z9F86hrsgXHT4NGc0YyRgGU
JZvpTimEtpthcQAPn/65a00hZzOT5BQ0eYZo6O+Q4QXOtj0gmmKlJekdpPSbC6e95i2G74jQ9dTe
906jrLn1jugu7YqhTS1JWtJ14rtg16Aoi9k4hfDVWCRHfSqTKRO/22LEvzLaHkMAG5twOozYCLFN
pXiPbH1BlMalGBIfWm3d/LOrWW2CFECoedJI8YxGhaDkMGCQGiGwYUzxot1klgqVzxVD8xoajhl6
oSnLIUKtW1TEUCnVJKkxhPUSQDFJqR7cXQZP3aWPsGCMDvlUT/fsyxHBwvgaVvLsqfLSO+NXHwpf
u1dnBa7vlxCpHvVMR6X6pQLrtmVXisfPruNYyu9PSjsWwEc45HiyEa3Wu0oai8x1GcDbxNcdUHvL
K/DBiqpETR5OHwKzDFuXUkaMVC7Iu4YRQEUnPR8JLPndO1ETJAOGtcBKZOehs1/0WBu+2F8jO1QH
h7PZUjpQiBKFtlYorbpLfK6Tk2vQnFia9fkCOaQaxDmu4RsJ5v0mlS0PM7pQfEp3KyrCStcJRh3R
e8Piz682xSx3ti9uu7FdI8rJwb5yB/gHna1zn9SB9jZxsuhJRl7o33N1qhkJXJwlDPBpCuWgabXY
JXesjmvRSFLlSLsaadN+7/UGUT+jHxOSvgwyGcTS9nyPuvWn1gLvU4xupH979OlukVmwnYBsoYE0
gpaLpsE8zoxLelZ6nIENhitt8Tuv7nAlPSvHRxTLURFxzMcSA2WhPZLMVjbDw3QOfjbCZML1UrEP
iyj/zL73zcWn4CkxA6GYqvBy18n4w59XO5G6xIXqZoSFzUnU17qzQmj6EhjZDAJEH4e7zqx9tVZX
6fREo3VoZBKao03LNKK1EcEDtYNY3GEPHQITnBE9V0uT0Q5UiGSi++bm5tPQlFIEAjUkokihxpTd
mHCLa1w5MALUGb55waa8W7TBvUiYbEHuKd5RQ7fssQGVv/WuIkOgOgV4vn3wN6z0nVoerdCrKS0J
JzUYZEF+r4MxP6sokZuMNqwXfr5GJDHEQ6HKPtm5vFHsvghbdi0zT+KsgKilHdfKsVIGNurh2PtH
53+RAejLFVAt8qedRrRNB4+odXjK5roUjicKy/K+5vlIJ7R2NqSv5C6c1/7E7o+fBLdqx4NSK+Dv
sJzyTEX8Tv+awvNhkeR884H7uzf1XSKc+4IWJNGGrtClpekfNK1wkFcFqfRHMyWJADvixdomsSch
SqXGuy/eukoEtNlm5RjKy+IYU/TvVXW+ij8wZmydZEAqI+1Sfnv+ZeVzjS4VFSV32OTpLXo8LEaV
q3LW4Jj8ScTW+1OG7xKUzp0obWdz1i7L2rDu0U4oPbIK9CBGcKWo8fMBfSHvKy7JXWFrWuChndqk
z65qYB6IQvc/xVUrtKg1Zt0TLDWKLvUXDI8vKktcwDHl2pdl8COXDxNPJXL8TnvBj4jwGNqyiYmV
wb8zMeRB+4UK0PGkPgnxJ43nM49XCHMoPpvK65SXstzBBGGyNlcCVzOMryDtJyUUURhbfewuBAW8
qhcKcYp5XXEjjZ6w1n6uHwYUuiD8RXN7QFWZ7MBS0LlzyxQlCp1odtE6jOliPSLNDHakDPvdq03v
DWZSzX0axKiggqsqa5jTGJybYeIJUlEgXKI/2EPrUH+x0vLBJNBxF8jQb9Gh69+cDJK29OK1yLXo
rjP5S45r5aljI7Uf+tsQJVkfamN7W+We76Rzt98mTGTRS+JbWLcodhAmh4DhoojqWWg4DLseSEle
YaHu4YX1NbsO9vx/JY/h76QSUTLiqiTN3vsABA22c22+Tp31aVWo+BocrOUnWPQ0mWgz2lvU9pkz
F2ZnFQ0UsuCsQ32ZGwhjCVF3nw25ozWVr/OqKyCv7VDJepDVS/2wBP3pLT9s9ZLzHNlu7RVLeS0I
1lsjY6QdTPOXX4wJJtXBGvCvkP83UFzk8VjTsbwP8kmh/xewPQe43c1/UysyTGWEGupQ7PvzWeDP
ATqPA6LWO6yb7GaQykmRwg+4olT1Z52pldiC201rZsTJXH4/+Z4aFRUa39VC4SSDUYGQoPLCsIFK
DgCMaNT5GusqiWZ5APXdQR9prMiPCGjUKQ4xxhm9ukCBGuL3F+0JdxAO2zdxJEOgWW50kAC+RKw7
656xgg/wOwOJPaUdb88qgzDql7R/xHlsjGKimgJ1WUMAkLl0KmDPPX4MidG8XCVfRDH1f+nbpPge
ib6KzNGw48OUUF5dQ42GcBwy0vCHXf6FqhGK1ldQMT3hOSa5DNjaXYTwjt7t9vxN37pQQyqKYkWM
mAGCkz4VQm8uiTXNoaoxWg4SdG2hQj4w85nJDP3XCItItKa3BKEEPkTpUQNvOxnrs1Y5DP+8kEwb
TbWFWdp4G+gQgdlVmZ/7RCFz8/bt7SAcfbeV86+uRGKv1GlN2z8+1dOPI0WApJyzoGRl8zCiTH+j
uOy53Hkpr/x1G6khAp1E3Y71KWQZU1bz9yEHoVTsu8WGvOFU+Z6ijJRN9hjL2qKyKi7Oq17BBUES
rJ97RNQfUXB1pV53dQeLHRXnn3VOUXYlBcXIDhFeEZuA17SUFCV4ln8XVG2HKjEF68rnRxQDowN0
b8xl7yh0KtRMg7G4CNjlAMwsWJZyOgMiH/dMOPr9kJUtkAqdMGdUoR8iJHJN+w+C8tMC/F3bwob6
DAxwu12LPgtmcDBpLZYLvWYVdCCkUYGrF0JpUV5Hb8eftoY9EkRLuN9kqVtVjdaytN+HmpsF3yDO
1ev2hzOp3oh30fSd2yhlfIYrzQ3uwf32YEO0dFDABeMWcKg86RT1iRm5J1LRQzGPEdDrMqdNNwiZ
ZhDbe5rfwmbAfjkYjC09iNh5V7fnT1EXFDdqR3vRmOlBcJsAbLl0Qn82267uMejJIs1LlsYAp2aJ
xrcPCcH4gZ2KMd3VpBAhFP6xEYS4Qtr2dvCfM/07MH5EzPZITrp3QijZw57+aaFn5+MJQbjMPo/r
iTh1mYyuq6Mungxne7kZXmc99gl1xarUT5BNn5aJZd70kk+T/tWyQ2xK5p7zIyncRCokjkHisSxo
UYyN499aMIu6rFZ260j+Ek5vssZcc0rIMQm8mL889PbhAvBXK4sO0Jrs0olDAB5/0OvPwFzQ45at
/0Fp0kp3sSxt6h5M+uuCHgqzaveMxpOF5Fs5hJ+RmzzWO8eVIUxIXgaeZnukcHVQDhqQyQQjVeaO
HObWEkNYWPXweouD5dO7EIGnGjdIeEVatuyDj7HnjxnhIfeb5vuzDsA1KiZu5etlcInvSyjPgOR2
v4vQ0JBbx9mOIbcGQPfdCh9wcBrJoloxrssPz9JZmcWwYYnI1W08dY4kAfSXZvhp4wjC6uNcKuHQ
Yk6dZB8tUOWdii/vNtDMqckcVlkAe53JIsfPNVd0qIbpkMStdBJs9teRhg3SBW2OqmOAozqgsPAl
xRi0slI9Wkf9w9FuSZ8Dn0zGxxDE4y8ss934xVdYFNYiD29Lukp5kaytJ9C5jib6IEACyOefhI1j
TXeGbVNo2KARu5gNzzMyxyRSL0vBNCR47/PtHWRrFBLy8NUU8g8y9B77MwkWX+Az4cPRlmkIhObn
0q9ovqbwdxTKJ2qhwqZ7gA/N4cSCILNwAxwEIWpxFg1Sw8U3AHot8GJKtIfUxNpVOcddbh7Yq55a
Fpmsx14cs3Q62T0l5KoXDyWwwRQjuCn2G4TODM4QjxMS7a4vthZjZJw9dT399LqJ3MmZl4A+QUva
qmwexVPnLrKpHgs7/TAca3Il35/8Pe8dv2kozl6zkl5GUpdoQaNr6y9QZKqKR/0Uv0nDFyz4ZHCC
M0e7aSYS86j7GL2DO3Dt1KKCEqXXfWt8GBRC8K4AFRNrSnB9fnaYCDXaBHtWO7y5wAEuGkDh7CgX
lEpUCI8BDbzHNQGkyEDjSxwh3DAIkiEonNg+eng8SRpgtijztaJUe0+Mm8mSuAK0qs6RqMXmz09e
2g7EtuKjvyNL2xiVzi6juTMzRr0C4LIStGCVcYWQNNNq4gaVwuljtoInXGViRwvQvxOL0QDt5B8u
unjTi1XUt7x/ovVU+NijMOaHkzLde0moCukncbQNhsT1zErKsTsHiz90U/AkQEie4QCqFKXTwDLF
bGi2EMGnHQb33QAf6BmKaIgFFXed901QLhNaLuHI1Z4O5nq4YhqYdNLOsTHlBMcXEU4nESuQucQD
xmFoIucEhV1nk1yxB/Hts08OMQMHctNKXy/LjGy0g7vhJHPv2r2TdktdytwPRqLRxVHjUIhj8ijc
z6fMGdVLPTDgWZjppqIWQpJiwE2iJVmRHIQl5OgxXty6tW5q6PkhwTlY4p/a1T/krPdkaUSIC2yi
6Ngb0l6joDsVg+LPdH9xmZ2lYvMeuvjLmwYQ8U+tIerHkC42/x8FbEuOA8+SsNUsxVRY71VsbFhr
D1aJwXwxIdqUt1IRK47TPTKLFfRIJBSxn1VWjekaGFgo3wSx0+f4ueWjNl4xievIyhP0JaBYteeS
2x7SvkXY1qYpveDsLUTXce8K5zis0iRIhjjfUuvMhJeKUZPC27QCs3SmxLtbpF909zpNgC114HCe
7Wp/BB4aicY8cjCweuLfBCrkir8HldIIT1YWZOigsoGCyjTo8ksal+JFZFSGihmn/VLAu/ZJKXnW
iya0WpbE7hg+2rD6fZ4o5H8eyicFuBnJkRh9EZPQIHbMm6pEAhqmY6argEsvMU/X+2ZKsP90Qd2S
WQozTNJopM9/NpfiBHYfUKSGfZkmy1o2jJT0xT6bESA65hyk0Ko98MdSNp+4Tam8J9nhJDi0ieUX
Rzy3eA7Tl6TAv46DoVFsXabK3O/haCKtiQyAXHroQdj0Mty5m9wC/iyiWPBHru0WZ6//Lj1hBcC8
GqS5yFkReoGSH618L0SHtekM6j72DCWInug0zFJ+JrCm3ngvNRJC+YejawCsqYYrSSrOW80b4W9T
fBtnbtrhkZLhvAovxMp35RRS1v5LPSaB3SciS72jZRFW1+dUA/dp23LXpgCoxiADI4xlJH1ZsdD1
IS6OGuugJvRom/MFyHMsJHhGnB3a6nhRMCHWkgK4+O7WP46RlirDVT8jQsSXrWLKxIo5A14sMz8l
NgqFQZX7ICsEwtpS1vOaiw7gVJzEhKqL2Or2TBcZVWcLEXN0jzvjazGmYSsen96MkNLEz65nkDux
1fdC0T0GKrI66xmChWuLwGalGB0iGgy0rEtmzqkSCirwJ0O/lhTz+XmbwqfY5v5ztq0lpwQ9joqH
awLSTdv9SvZk4xolp1Xb2J5NXZtbbc0aHnCL00r6oG05f7DxLQxpBxLFtrB5Rw9GZxWYKP8OgvPb
ye7swC20ZTneLH/vwn9KoU3G9mfdpkd4uGKIVY97nFMxLxbUmqzh8/IUbIqM9CxgUysKfVPHkKku
kTfIrA4GNBLhUz4q2h3/lWmai1WmtvxiaEBR4SzKuEkQvUdYqxupweqFvzzVnRWS+buk3eY56Eap
EPI//FxjPvfLFhkk8sazN2XRL1uD5DyXOSZQAD9GIfgGlOFTnhKtkctmu1hbXwOG5Q5in04u/8uC
OIHI5C2ft+udx6U9mmQ/TGRpGfzsOTg/BrF5b3bNqyEgBez+D/Ldn6zS/+VZSZO9kfQfyBh92AIE
6qpIDyaAN7ASEFcq98DRyHbsiu2zwLLUGcPt6XrDdRU8Fczg7LSvaRaOqh/jchPRGNnyHaGac+LP
qjwlAhPphULJH6QfPrp6vmY1GwVK7crYvkxZtRW4rUHAg3qB615EhfFiHTHl/cvDqTYCpauQIpXO
H402yv/I2SPbZlegBKinD8BzX146CQ3/NlTHd/ZASznZeStMYhPz5jiW0NZSOBAu/JzeCfWPw/M6
S+6gRgMc0A3aTTtGG08RDmu9Egnsgc2lRE5cUWYzbnbq0UeeAakego1yBi+HKy9m4ie9Y0q2n0pJ
qCYHldthbxMR5O7XV7X+gxE4bEEXci26x8nKf58paVxCobSouJgqlnCXL5Fs+C/Ld5zPJ6bjfv8m
5FECPnHQ68vYYtqG0AAF5LD6CYXFL6zgzymaAOOe446ivCSpNvWpxx9IxnScBglQr2NUVhHZYGfL
ZYr/6CCM+005zzeGFqLkemhnBR1ys0AXktlw7r5O0q08GIef5zCdhKNUGIjC47nWN8CTBlW7Fcz/
lEz05P4hZ3P5zwyTs36J+eW7sH0JWOwNhQRv1RWTMHrIaYYQGZkxQTpDoQCFXi1hfL72b7qCm8o7
Isgf4WZExNiug8RAk0jCSWoStL56ExEwDFqC7iqptg3oJPiXgNLnIvUBVvRqEoruYYPrJxu0mJpF
ELW7wKDWP2vc0wUcWnyP3teSCNa82RyzJNmlnN6RsCMR9yhGLtvAA/0nMZ5wGD+hJ2pPd2n2+dGT
wxNlTA2HrqEgiz9vOUEZBcpZGqfb9uFsGyl57sZFr7Mev3iE+IK/dDhOc2VcIma+1a1cUZJM9pgm
v2w8+qscxtObXK3u5g7Y6D65ZUu9p13207TeCzQfiFgeHXF8B93UryvSfmP6fPNskLnYHByZL/Td
ODBATlBx/t+/9RvRhBUxTlE0/zpNkrVrwMbZiYSo1dIGFiIZJigOLCdsmKy9iolTUkauEy+RI4q0
QzKJ9q8DR8hPPhBOgfePI+N0AFRN0C8osoNO4zaaXZxJHPhvwk1oyfQi15ZQ7gy5ErXuumqHq372
avagSbLZxwDKaoclM+5Uyaj7lLkp3gdNvQQxh85+TyZqTOV3IKzsDApHbFgOyY7gw2iNlB4mAqyy
twIsucUaLVOXTd81TqsCDbYrScEoRo2ITpDhh1gJ6COvueJD98DfSIZMd8jTml7uQRKorBN+6P/G
gGJJLCUkBLkiaaL1nUanQfeWITkeJUbUfvE3vhZx40btxCsZ5VujaWcUPnC32EO/98oMKorMksE6
zljbhLvHkemKZqFqexl4HFtyeFDfB71qcW8zxf397Len3vvDT+o2j8WLIzTvITiWU4O0+TS0Jt+M
IaB1erurQpEbsU2gX/m9FmLuBzqbvRZR9Q4EnfDZr8AfmExKAi+q2UdzspCxS4z2XTrrvNQnCBn1
Lgxb/2+8fWv8SvE3kDWIA0qH7TP3Re2Tw/0FeZrPe5whtLfcHuur8YY3x5gtDM9XKfP38dN4fo9S
pDoqu7oRxysW4w5etQidUC3LQ+gvnuuOxP6QZ0KJOpmtcw/6FqY+/g83u2t2qlkgFyBSrVP+zffL
sFoYwyXGn+frtAaH2k539B9vEzbAJgUJuFmDSpilsW282MVvdGsnaYrvTGBNRo33SZExBoR/tTLN
fvKDBWudPg6hZWV9TGfKpGk6kOCFBYVVSQBNlLRD//+I+uBw2vBUL9GScg8pkwECrI2WXu5Rs4Uc
20JceH4vL8ooXdIMWeEzqO6Sw7ftK/N60urBbXa0krA4PwTu4OH44ODhg8xPE3K622zbHODKrKRg
A977Ww3eEwM8WgQIR+oo1/QNYNLoAlnOxNhg7yEOs8TgWFqnCrJfH+lE5hK+Mx1404S5oFHmCMHW
jrUZEF/jyX8hWiCwvLw6HNDoC8CID0HwAsiyB36LuIDR6H4bWyQZHVlUQ2nSced0JryhSrcJua2q
7oE8ngVWUbKpwFTadYwV4Z9aKbg79g2V+4fCgUJFyKvkdGcDx6v6fhRbM+r6k5Ev2CH7WuknfnN6
HWQdx1BoEYu+FVIOkG8a3b+uWZOU88Hi9ebNtYhTToe7O+GBqdN+CzcEsm6j63n4GJH5Al8F85bL
WAjvojj9CxU5boX8rTQqQ54khGVmFS7yLw4X7oyNlil2xaefO0qne/bBXrBqi6z4PUDN0DUQbQEE
aS5ZEgzcI77LRQW2MjYHNyAvOapSsl8XNXZDDENd3e7CvLjP3n4B8ILzhynJavol1hCA+/D82cII
MJ21GwT1d4VsuTGHpc6X9/W6fvvW0cNdszcsWP2d5NkVllbqWWFdxpen9C1LReX0wX50WxdwTOZD
UDbvRGKpj/46aiTkw/uR3/Bsfdm/hJmeeyqJpmm5MNJAlpXU2/XVH7QelYJ9ADHFStUaix7/lAEI
MVGpICXvUoBoTSXZuBIv0LZ3vXXRL2iDCK/fNevyujOUAjn2rAQ3QLl2KgCVaaSaE6txB6vz+LCz
H2RRkjefkxpjcWpotMlSN25JAH359ArFwEu7buTZXd41voNQvxDofR1u+FtT3XrgpANKPh6fCVI+
wAJN3PxY5cWgcobPsOTzdvyj4fTrB++PXBC4SloUXrQYfkxU+Dt8DJE1VyLiJFB9lHvHmqDr0X1O
ocBuiJwkdk1LKRRsgtrXql9JcGk/tOR0oBVj3R8M56jPo0Q75N28MiHQgO+xviLOvNNpqpYtGM+Z
UDa1XjHFggp4S6KwDsg/o8INpvcvPEOLEsoI6HFCGe/eXbJM0ugfEWWrh2eIHUX1J2XxEcDQMKQc
W6FwKKS4a9b0H8jsUW0m/SZgW/ggShg0YlnoQ+8nt+mWxqI2Bx/rfyLIM7GNBfqCPYe0UBd4z0Hv
Xp8ifZt0UqMu2vv3ResoqkJbPTvQ0MnDXJpB10xGS0lV46OUuK31120fgLJKdj4LL8LoZad1rS7S
vvTa3ZsqymCwOz9NzUpIr7tT42kZ3rwPafcIC+163r07b5LgMSS0lFqq9TgpVpSImHDCsKRDqNbp
L4SvskEm6NPHS6oXzG96pktcudTvNlmtoPG1/54aUBspQ3i1n8z8nv8gJOl2S4ymIYW3UTuHOlBF
xmS5M3EazOduQG8vIZRiVyU4EJWJ3+J94MCRzDsJQlgj9yHuVY3K8KBeRD0tLsQDif97I1lLc13+
ud8t9jM0fnvUAtCI/A/9QqWDFqMvFlxNbVjuybDFchsnOQr++GlCs1Tp2pqReTsL0IbqucEFlUbJ
/q5+tarRMCXh92iFEsQUXXpSA+IFmGOJg7i4KK5FlN6hp4H7TQuaC9YB7Fqf4679ixx7qZsLXLDb
gRlqKZsocgvCcSGlFW3wcUFaTq36Ngm1yUXxs7bYKmtTeOr+0h5tc4IE63imPfEHZHOc30KJYzln
QGhak38DAb2NvWvlIs+u7Od2dji9Lp0PpWMBCe/y4X8ePCXGMFLH7D1unDrIff9UefbDJpuJ8raB
Dtb7tbtzY9LKEnt7dr7DItIZ/dnx3cMDcesVDtzZ1VSAZNDPmPJm28aD5BJSugaHF4oW4z8NrO8h
tj1iPgSWzPATMyVc3k/IVFKcXO9qF2Aug1oqQ4OsRWIRkmkQSnh1QHwSWE7O1L7fMpLQaIItETP/
Y/iizQuyF48pMIrUP85SgueHf8cFHaBi8bgKV/8SxIbW1kLcqmaDOzUDWgMwyAJZtOqm7VYEpYGD
6sI0fWcEFyt+yfDGrPHMFoiRkNIlQwY+7kxL4D1hBeso4dEnYUsciW++eJOXcRF5r1Fpgla/iRE4
syi0MxMEE8/lJxkcWDMTWPAorrpZFuxjPh0OnDv5GDvb30IvxI9HdK7wUJRTSLkhvpBrI9C9unug
hRGXrTH/saR8QycPU8kB3hARF8IIEXyMbieA5PiFgQx7Ic+2YaPbjcBJyXCSDny8H1c+tk3DMBj7
xw1NUqynTYrv/PtDZoo7wUl+6+3Ae/0g6AnBzv4LOpMg6KXhrIamq2fgh6npsU8Q+gPdVOuj6T2O
8KcV8hhKcKODVClUrif81FStR5R3JOQn416JbFQRPC0qfo9ETdPhGbQH+8xxAINVHf613Vln1LbN
AUIJV4oE5zkncn954ji4M3sNc4s4NYIXgykU0GXrdjecs0AMad9U7bwBZWqF5O+2Ecnq+GKxD+F/
hPrKBYL9X4KaE4gI7ohUKz9z7w0FuNlh7FuRXFqu5vTTrx9ULJraodiZ/pbSn5lP+zHsxXs7zrp0
k5kZy72EvIS+dRARNuSWXpPpWUh3p84oXmFpT/j6JhkS/QV4SsBaUsvlYDC5ag6K2jepr+7oIOrp
SV5j6YngX9LqBykHgmDiSShytVzxrxH2tAPU+vH5q7+qJiyNa2RECwNobX891DyUudxBuLxC9s7A
O8k1vUPi6N2M0rJ6MJE0H8B3Kh4X5GV8qQKI6JQCU7cFJCPuMgdrQudNhInyfoWTagXtC9y20PEh
Q87I6PeypF0c6k0irK4DaA86Qg/AUksHLtGUplDcMxSTyMsKjGL0Cc+DlKK8KRWu/biLVP/gl7W+
djEA8eSaQns+2QUMf7560C88ZE51ZPk9Zunm/5kEbatjRev58iZQB9QYp7eY6kUyQC/Zf+bUSUqb
Qq/vriHUW7Qls+sWjr/a3cvsjElEvgElE5bRLTD47Zdmo25LVSRyOtHOjCRxsx70UcKPuWe13Z7q
NfJsZo3b1s7u1S2P8x+UZKO9FlNuyRSjqBh8QHzfleaB66xXzqejQbnP4jHlQOr35j0MOCjS334i
uHpqD8yg405EkRfQZYP9U4Tuj61pse/njQR56WZZ2bb12jfZ8k10Jp2pmPSCYCIUs8aQjtVmNCVU
ZppfgLMpD6xzNwEDbz7i7BnJbd/Vji+exaF4Oo6Cb95ipUe7r2SGGt2a/ZCEs7j7bQxw6T9b6nJf
+WwS7Bth3kiaFskvT6WVuQ8vrnBs/f5uJGGnimR2feE+/wDQVpEa0lRBjMy/2cOmGGB4S99AiVen
2I5yqLUG1g4w/ntRzdC1sGv8oltYvEYnEuw4wEyJhpcEkJJtEBBzDcJWwcPV2Y9zZNAC6NRBvUHJ
Q5KzJmfZpIKDp65YlJ4IbxxXTZAha34N8eRY4mTkMFcYahYgEKeWwZyex/brcA+EsIwy4ZKMD77r
vexf4JhPwa5ZhUGoYFDJy/MxQ1mbhqn47wE/Xi8bSijl9LWlG82PYOopRta2f71ROascMkRQttJH
QK+3gHn6QUk0int0FYPgstzaRIwiMs7pS5bD03KLQnAy91ejCAx3LVmT7h7xGV70niakYJ8bZtyH
ygQXK1TssqwyCcg3ep6BoBPfdUq7/rSvOyEzcbOYMhYYVAL6qcPnc5wWIHgfY6tRoIjC6VoUqAs7
kVhcv7Bkn+hy7xA39C4XuWf8iyJBgPSnuVD8rN9QBsP+GWGOC6UYixEN6hkyPCn526WxgBePA0ek
CGLbzxcPCc1tXB+FAtI0w5CzpHJyY/Okm8qA2cxZObYMcm6kmHK+MjVqclZrKF3Wa7RwIQJnVxAq
0cm3+srNJvoIo3W3xA67zoGmgiRBatVyVQcwtKKEYJRfIejBwEMiw3M29meYcK5TxPWqoMU5Sv5k
RrXwFPLX3fjMjgX0pyrJM4p7Ino1LDjQ7L4a8A8f0DACSeoQaEnmOA2E7DMDw1YDSlKtUACMUmad
m4ki2SwcW4CFTnrVC3TooPlK5E2hJSPciuuhgMCAY1HrvZxrUO8pDzXxePkdXvr0JGaSxEe2HzFp
laJ98o1EsI8uYvaUUvru/0vnIH+kaLvIVpf+Uc/Z9ZqALMKEWn4+XmHa2WOnmopDQCcQOwpgYkIE
O1HRJyXD/6Fe+04XESrlNs0PJMEdQvay05aUVaR1ljC2xGqoMkRL2ahPX8H2/WjoMCKgxMN9nN0a
+uyMOEI2tYAvbTFcA9pLCcZbXNXc1hW2z3md65NzTuK8+P4976Aqm0/A0Cz/37vEQtLotiCxRMm3
o7POSKHi3aD1v+uBWP4B+/E8G7aF9JCYpHtdecHhkjn5G6BU+wIpFib5BFlO0uMf2ZgQlnPSIVw6
W3rT/d7sTJmhzwWFd+23mWPNE6LgA1xqrFvTP70ez7xZES9GlYCYWT/9COVxfxA7yeoJgwOWHnqr
NiXyMvIx/SNjtQJxg0PVxvalCzrXitApdrxkWjAL5plmrPZBgFjkrLYRfTCOm3jbpySo5O+b726Z
lzv3DdusWVygkqZAnuI26KceYzDMny2r/r5gH26ncLZhk0hg678l4j3PfZmUy2brG+mGQzjKkGoh
hyHpXPcpP637SHVzY47AoLkj8gTsgR17ci3kVhF5dwSXUtMI9pfxPQ9Fn1vAFnVqmR9144+7sqJt
G+P7mnt/Pa+LbW75pvCEQ4bNWu1OiP5BLVcdutc8PnI5ygmfO1EYVJ7smooRWgJC1sxBwjYIEvs2
AUSE/mHnz6jrUdALFEVNhymgI21M3lFtuRCzDyMus3o1B3API6IvRxf1e9M/xGyeov+Mydd5phZB
KjJ8I1SthlJ3uwN7jvyvDB5HbqEY5BP4KXb4xlVSv8mB2mYbBytA33WEN/eSrOCahfwT5W+edlUy
gCG65hZT9X+N5J0RuMTNIFwjnlz1naDoVOsSUuY2Ic/TSeAxib5+DNw8Y6WsA9zbPi2z7PxjIA9Y
atUbnUbN0zqlEBeZWiuaD0koVZ5l3kfE6Tjk8XC2uneG0GU5Hh8YwXFtejzFAtQAhgp5O/bKU/Nd
tK3NX9n/JPfyCnm/W5Pujrz6UGbGqENA8RGzA26+wo9AC+hkku/lKg/WifLxgzBiRcokRg2oQO9X
I4LbhTXHGgC8EgonG7zrCIjsHN52+gWOPTJrW3fhMxpCDC/zkGreAih/2T0MquAV+CEfOjtnujZl
JFciZyHMXp6f4tfWEJ28PPcEycmhcmQq26nDsMotLiYjIPFszFzgeir3+C6R8r4ykZ1YvvieH3td
39gvjkQXbiFSTemV4QfdY9keGHv8+pvBDhVG8uPD//S7zD8AAIB/3OlP1K2sqVU8vJw3q42TVt5p
OX812gdYpoZA3keDtPRS1US68pf6c7DdlBdxWaXTYOMPi/PPhj91it4H7v+OZGQa4dOPZvoZ4Ys+
qWZXv185XPpCoxb+NZ2/T3qcSuS6+qD1pvZSe71+80E4NqIW3erUMQt13oIQHQ+29nJKZrOMwTLu
VlZGMQYYSSlQA3q/SMSR583+ERvduye8TI2+AYUXZ7rOCsD3MnojKNlN50PdGbNN3nur5OVqJgHi
r7NFZcmOdh9JP2EG0iPl5WjyJk2t9wr/EbKSKZBiFkwaoG/JXYvGavzRZb6VUEcMUce8HkizPR5D
nT4yNU62anb0HtCzQH9H0jwJMf2MMqI4oSq8jnoKxwvxK01IC1L6n7YE5VVkDxUp7X9ut6k5ejzi
IMoYYgVe6YF43JWDFC1SKdwNEV413saey2skOfclNRpAcTIX9HvezOlGeZowEZpldu2w5xqo7hqE
Xf+ea+2e6Y2E/LBAscVMSt/vrcDKeJs06l1woepTtQrBFeS40V8TzvvkweHd6vVq8HpYcFQRfElx
pesubCLRFSkZnAidhm4lK4XXqcMqVhbHFI53++DEGZ3QbfGBFF2xLx0eQoLcv6Sa8CuzULIWpT7N
d3C1lhlQJIiZGKUdDrK562AzfehOiS1I8OZmD/YU9EFyX9KUDCXvmfNJis9VaYw0wTFPxWUl59+k
PTuS9qXIQP3CvoQOUpMpjm7uRPCV9GDHmcA2Z3dbtlzecSOR7sG0sX5mA6CAO6ETjRsUfH4SfFn+
fHBtpc9hEw6Gb6c1kcG1vEbqsJyvVfI1Q6QI6fcaKiR2BYfaKpGF8XPFUmiY4awKqDo7jQ/aDtQY
E/DiacODyLeJiqH8jaBsRavZEa0SiYpgKeV8QyYzWaOrByQdIe5i7Jv2QeqX8mqPJQXKowoppBmX
MWNO9JKuHQh0t8VjsJzLz7tSsm5dOCbLkXr3OHsjLykIw1TnOL1vTB72MVVSJB7o41EA2onImrUA
XREEnpUOj5/NF8XStrCWRV1DIaca6smGSuTIefqUY63rrS+jOHLEUzAxYXId0urOaih9sidMmbFF
S6ZPLy5MHBXnMTDrdFnux3YiDYZTzEdYjYkm2XbtFEQWYwBXwKOYjc8DYiJKxriL3geUAVes3pfO
zxCCiRAi/G63xCQKqmzQPpyuR+L2Y9dxZxmXYZKZ3LYphWdynZ/uhCflFl/1WV7WdkETgDWzx8Wn
Zg0WdWhvpVD35FS84g+1k0UYeG3Bl9Y7TaDdwKPVBjs8WjA1qVDSlG7upd/LVYyLkHhS1bp1qQ1q
CCvXGsgGch9pM43fpcveu7svlXa9yI6ZeTnx5q2KVOfLiQsmdRwot0EwT30vB9Ta55ISdnJgOwuP
cQWIi7A36k4FgBqN6N5UwuAbvryAhtH8QCVLXHuV7Ob0dG5ZuQBg5cOuasAVSnCpd0p3CApiKn8e
RS/8R4980I+1nOBXGWjCdCL0pUyyMQA0tvqDpYD0CnFOVJ7dh60JlkSgsCm/dSXd3bwtvdjLB3if
NUtIDEIOx7uGK6A+1dIptwZCjeWoGoRMQQ5ESGTbHPO74PbhtLdc+Njod+S8QVEMJYLeTKwRKb/g
ioLS8u/JWkNvKCvCZOmLs8eIZ8gnyUFXvDHEdaL2htrSn3lLWDgWno3VamqOpFsjRrnZS7xWZ1i1
HAB6QxZzKVnCMsPyMejNdN/O9CH2orLLliKuV8sru1zrMtvks5r9dbZEKWVyHKA6Pmq22KCZOr+5
l2xiBgJfGEGel+ToMBjgmOKYB4UFvlWBT8e+xsfKw+CIoBbbQMh52FC56cnWawgzEG6Vn/cy4e7G
ZNEqjuxPOI9Rz5MaZb332AowXjtzM65ywKInmAgTXOMuiJl4rFd3E8lkReVtxts1l9OVd9PKW6JO
WZnsgX4lYfeoFEynRMXOcrpSss7ADxjG29p3b1YCoJk+N7hWRr4zDoELwnjRnUsk7ofxiVjwKOzG
8DmpKhdJKSg43d55vVGrPQ4b6IFaAGuH1JfwQiiuOhBUbRxE5zfpuCAWHwx9Hv+YSrbuxVpBtsgq
HiKB+Ftq4+iQ1J3LOFhFr6F0W7KIYFE1SNFEYyBgyXNfBV4imi1L+JBP4IhLIdcoxdOCWzHzaQKY
PcVkFsVSWTZZq/cH3STQhh87RTc6Ut11HZllBDYn8q4ooou3VyP1aYTh8KpdSxDTqnhoA+HBWnfU
iMVC/yThlewN5nWaijo8xDJ8iIL2F1/tHR7Z/mWCYY6yiFFCdyg5+/NzLxv1cW8QStzcJzhQrEpN
97u/L97o3mh/op+eaa4e7RoMdMjVn0naIX4HJI5XiNAyppq/AAu/K1gYZTM5wxxuUKgMXAoWDlZm
SWClY4iKl/OQtYnVy+eOTMcVwM1qQ4E6YPQaNz+9gO4ICxdT9j5eiXfZWHF46qbivxX8jB9i/CqY
AcAMqip2TJ5iaYr4Dk7OQ9qia296JI+B6azYiuoB46I6WfHXSDxkb2WAA12o0UEa8YxJb1RY0iMx
WEip5Zxo/VrBzX0T8GZ4zmGMfrcEkL6meiEFtdjbSW952of1TXjaX8GpTB1MDdfX9wFotey0Nv9F
9AU+xbiudg43gvGixE/QzXxnrhBRTUPCM+/WVuBRYeW5VmHi2R6w/g2NJPyf3KuhAFePUm3nIjaW
L5X7YSphHx9Uj3BbzGyvA7EQtc9i8ylIuqTUfo8ximzzAudDJb4FrDweHhr60Nut3FQHTetOA8oP
XviqbnBouFJiRHH3EQ7rqtdtTC4zGTxBkDA70z5tFmvNHgvHJZGf8/CDw/vQ4cz9o163RF5MsnKo
OL9z8KIFyzuW/32SIAFHdzCRM2/OUScFEnmpbglUqNiYWwoGx5diPPbIINy+iJXD3wiRcMHGapM2
EwhWfu49/gwvOD/1sWnBMUSYvh72WwD6BtR5YQ6q/cwZcYVhqH8UO1AecC3GoAcqzYXiBOiTEklD
sNF4FeSZ8uqHJcvGUC/Ie0WEpDSEuosUe0k972buWjZfVYrEv4+zpZKKtWVyfwIgSXawsCu/hwpx
4CARQDMAIHTe7F62G8lUEyjrz5wPE2R5C0C0S7vcLdnDKeoT7GBgReC3n65kLWUuDYZMMzCN4I3I
BP0cOO1UO+l7UdG4OzL/8GjWnoQ/4E/F/N9FgJDSw2u9EwL2xptRrAdmu33mjkSKQu9ekyOwr7/i
cEhK97PiuUgAiRdbmmKOB4V/iU5Txqedt0VVOd9gSliUAWuH6TKgDTdE26s9VSL0XvcyJGAIQrOs
cbUd6Rnfr+uLLEjLuYHwvlFCQhQPsngXk5FSR/BdDaGpgGJ6uy5l+e8fVNqHQsRsWjngDfzUo5CD
0WhpRt5XVm3Iw5Lvsovt3w9I98SzvEpUWsMZBlMKWogN7AkSWcrksKf7paV338dmZSnMlYYKW9ih
hvD18YwCzusTXtqeI/qhRH1DRhePH2BJ/cKRwIS4B2tpCPPNXFtWW1RRpCJH2cE4Xq8me9dj9ZdE
MSejqjQOTfkiT9xmUQdgi8ffmTLi8YmfE8TxCw+Sw9iL4uT14DyUMwnl1pnZiOt5NzwJGjX1eatN
D4f+j0GuKnWgvS4NzYUuAPumC3WtbcEXV3T3WJ6y7RYBWTSapcrK+U/F0IzF+CIYtjsprD/fm2ci
7YdhoCnNB/nQZCXcpdTnA1SBMD9yEFV03vhLINh9gE1JEuERk0FlI7pxo/SfCgqfDuebyZz/4Zog
BC1/4czYm0tMlHdiDdh5adrCJDrcfWyIrqyQXDetCyw0/6gm06+glplnId7QmrufgkpRlXz1mwEG
zFgo4Wpt1H1UWgmKrEgvJCdj+NLrXNSxNkcX+R5mHry5qSJmbXJwuQCf5mqoI5QkVEuoaT4H3YaG
tTVoOYpgep0dadm7BLbSxlRmfGAQ0v75njHwSILwUwQS0+joGJcLhYOiSRjtuNQNiS1Tl687FRhg
ZhO1NQTIy5b49Z6MRPWZv3ocbmPNtCkI/La52BBAaSEIOnaRU23vcyICDU+ol3iMhd74OeBbADDp
igTcDEsT/RWzfApPZfOpt/jcWT/DIOjcbLaUpgAmHunJsig1G7mvgwHcjRfYCuDiwkUtnwpl1gft
3IF1wlJrIVvvcEimFjTCBsYtfAjKlhPGbrOze2DF1Ys60FnBcl6icugr5/73mVI/V/W9Y0k+DmbE
Sv+d8CCtkZ91aplEdrcy3j2A5ff9pjCJHDJ3kynOYdNNCh01ad2AS3N0cMghsfSx9PK2q4e5gnaJ
mVQf09WasQ3xzLU957OJ2gcBO3KbXUH4Z1aVXvMQlp3dqzKV7DkL+N3NukbxlQAc9R8kK0Y9KmjR
yzBOdwfMU5uVMjdc+nDu9v5/IuHd+tsKRUehF1hbVG4DCNZrik4FSfdWFkSG6H753jAmA/B6wmrf
dbCpTbZCjcpkuRcIO9zqsV3KrtRy+xy4W3ewSC2ye5pWZJ2xrKCuFUhCuZ5x1qpfM4Qv5LPte3tZ
rOY/vBLOMMFd4xvo357TX6hZHcuFjrSU3BrSfedibsCL7eJsD0cYM/R3/eqP0RRcE7+OxKPUKrSL
n1G4NqFWVRoC2ub6ol9HX0MsZ8pu+BNJ3hFLcyIDsb8+DBK3xNZkE4D5GThUNi//xPHwUR43hlb1
3IINfWYKE7MfzgVJM8X718K9GdRYB+10AFlfxpTIpdJud5n0M/dyMWv+2mrCuRE4WYOdadsmA41y
KzS8BLjQBk5uze0ePlvABzWmmCj/1bBlAyiGcNo83yYwPQzMf71XCH3X87RGGvcfMYS1otBJzqDm
Z1m7PAXbBeH3cKKrYVRriY2l+bZZRxDSt+lUvLT5dtlFhD02ibpm3Z1fOzp+2lxBrpoxys4G58my
Y3h6yzvNUXGs1uv1F6oc7YyrRCNwrkEGIFnOasXH6eKPSR7F0mDDmWFXUof7syiFmEzUHvaoM+B0
PzRiJpOCdtUzXcsQmu+y1SSzZUb0zyuc62RaZzaitA4QBIja8wuDB7q3woCHPYgta+jzJQ7TNSh0
D6P9avyGWD6AuDXH/Qb1FX1PXiWs6jQ+CAi4kEuMAYQ2kvoaPl3KEIAAebMq5q2s54yqDuRJDNv/
oIh97oGdywupPsTSgvieFVs2eZIJM1ikkOR6s8fwOARpL1gdkXXmsfgOZfczdRN1+PcyI4/UdcO7
CkaWZIEaojITd73jHVWL5vG/e8cZN8m+lyP8DjgThgMlOKyBnF/2De5BDIy9NP1qOp08ZGL63vY5
M0qEDUkG8p3iia/ljUvPN2aEJBVuZphmdFO8owtQ98KR/OUj6gyN8f8ToJ2jI4HQvasnjWEIPTEP
46PnEWfn48lPYrogzSW9S9V2/iSP3heKDkjUgbpmiOROuF8wBtpO+fgKnfPkx0Lbxzh2WtBL56ST
9r07W5ISg8pqB0yMw62U0VOq3mBgUiIbvul8cBOGubN6pNE5phFLSQTt2tUJdGIoysUSIDSjpFsa
hUKnzDtAxPwmZlwKxm/NysqjNfPxt3axnqKxAkWLmEjJkhUQE0f6vVUfwTqH4y11p3e9al9UK1nA
XL7AoZUMKW/846Q4eDDlIg3lDBpBPCuol0O+4vYuzXRw3PTmPgLtddswJyfK2zifcQbEZvKj3/2a
RjYdUayZ9m8EjHvwrKswthbEnlrHnybUveZvn4cYgA8LExIOUQ4Y9JwsCDRucm7QGcVo5GoAAtjM
lxi7QGzuSnNGuJ4SiePbfN1BmVGEK75Z+LAzuqb7069pwM2XtcUYYSvc6u7icegWULfubl6cxNT9
pOjoYALqjPfSeVrmoTZmh0NuzuLmUuLGPOtpM0y+oXRQQt1FyiUz9UauGMNZqmcsWAybMi/IW6Mi
4iprnfV/uds6ZjDSXqEH2xJNY8bP3Ti9HJ6SAERgm2yqPlL1wKEmy9U2LN7zZK90zNsFzpcrmZ7x
GK0x2n3mGkW2vRpXMCSo4ABDmlYFAhZlxIBC/NKuGT0QLT8CX/bAzDhE9v65wod9u3iqzN8VTn04
cXk/J7+XNML1uDeLiZFmcqm3CJITMMr8ypYjAlhUb8/4rOqrSZn8c5tmRZumj+F2unvPLxy1OHXA
DekO6M5TDWjWbYOrNTieC4Bq+1WEjqIvnVQlG7JGNt0AJLanL9D45IsauomNSYBGafxQBQQHtXNV
aT0rnc++YmebUfN4nAyOC6dQRxMw0M/NX2ws30CpAHqh6NhYPLnj/ZQbHauV/xTstSiQ4QKjf4Zh
jGf4s39egJiC2BrraEbfIWTmE6kWA2DCoaqTalpQ8/19Bu1uiOI5NdTwVZbww9CKUm/4tK/l3gFz
r/dNom4j0pbM5dZLxI/2fO9vP/VZTTlwHNU35HlL5J2dnLZKZfjhEK5uaCEck3MOHzcSUqYIoT3+
6ijrK8bK3fCsMj8mFpBROG3UVGRTy6lFZbAiUS/KSaYlTHISARpNjzpLRVpVEhfPNJMs9JJ1o/Rb
rkv4ZbG+9Y8d+B/A4wCW+b3ECstiNBXd+heuTNu2jdTc8LU4pkpN+5JqbsM3S0a65dmwLNBpwPmw
Tu6YJHzjoTRXgKHSQcbMrMfGFU0oOvlZTownP0kDF7oF4fhFLC3WsUjFzJL8mP5UjsBg3rLUzsfG
k9N53jmtIxCWfi0iqvBiwuQYnjCJbvkS1h52oLoKae60frB8wZeog1GRiDRxZSh1Xw3l9fUGRG2M
RJeCKnIQ+iJjJhl8RDnMCoTg8058GWzJ1xU3l/PHlReCb+vPwG4V3a1YL9v3/kWFVtLJ8r5KhS7e
b78qFg9xF3MsFzXjXqDiPv7pVZqyCtIOCny+RVMSegrY/0z2UEChYfm3kQyjI/T+KYdiTqJOmKdO
AV9yCxCdNzsZTOwJfrhTJJyh8y0sZf918CfcZ4kIv/I+HOIuGljsWZeqRjH4WKNOJmxXbvH2LFXt
rOhnSXTzadulW6pcpWG27w7QX/stnYHci+7OndJWsW+GV1Q+DYbqKAnOqy+5LDDTR8iJ0L3fOBEM
A2KYDExmIIqRCy3mtV9VIyZvUFc9giDS+XhAGpHLaUdOyAxbNN8vq7vT1yh6LuNt5Cdd2nDt8D5A
LEpS0QNkvuTzKmQUlSg7w4sg6XM4QrLHHjUwtoJEbF2Qzb+GwqaodaDzFNEmUEpyKuIMQoLicAJ0
JyRWTClnZpxnbklLb97VzttMLD1VSu+H1bUSFgt81igd34+r4MWY8E3/COfsUS0FNwCC4jZIQh5i
HhIkSCiSjEmPx5sY4Mlcns5Qg7gPFDvuHVbSwC8/FPUfRfFmy1JNz5+ioWu1Pv2y5xEHCCjTEC1z
rYAoWYwFFlNPf84UqG6bA0/2sinj/6F8PicxuzStD2TnuTmaEaXqc1PoBFmZ8T2XkXfSZp3XtQfc
KKvfNax8VZMv8LXZLZz572LbTk/myYa9kLrkTqBSW0u03crxlJfm/BmPXeM6oVIHMrCgucX+Gd45
M5bmjkKPRV1U5xwDWQ5BUZIUsBnYdo8IyYY1M5k1R9ahd1Lcq41kKlA44fJgLkLgIMlWgKHDms/X
xI5ygsaApsAW/Wd24ho9Y8u1iQqmuT2YxxjsP6EuaT4KZl37otC2UyNmRkojDD3AspewE/aquYIC
fVoVtJANHI7Uf38+6g8zSNPm6DWWBeOZmkHE2n1v5YSiyHy/ySMIoosNbajpc8RAZiWjj9UtI5bw
LFQm+MouA0Bnws6uMnCUwDwCBj8ED52gJcjQ5shuEwdth0XLNX/8eytdHy0iGtWSd4DQ+m4XscjU
a27bnNmOvxzwFWBBmpAD2VvS4lOXXZxh3kChzo8Q4aHpkQhJgeOmIJZGgfausYOPaMLNWJrvrnXB
g9tsVJvzkmIr8qJzivOYbmxpT11Zr8o2dfCgtATD6XR140TQWCiNqqBuzil8ksHorz3VYLSqfZfX
3hs66PPG843UUbB25HLY2LS0UFkpHArZRNRGCBO1hUtgRP2aHevkSUqtQfqYeKLnbOJv4DAzA4R7
A1/Iv08zRasXfDEM59YmlJW4LKfBExN1Tzg6yECrTgXqDoZSf+Cx/2LcQUVE22qpvk04MRinWSBU
WncJfejuJzi/Ts5E4Knsmn4sEMrEwfmfIYFpQfp1IFkv3vXltfF7qK8CJGNWnPYRcWR3ldCXh+AT
dqpgooDMSYGKd28nsxFaeGkTDJzwwLSjUNr/Rty5mRTFSleDFpFGxGrn1p7eEqm0GZIRcU0SPwaz
n0J73X/UeeXMX64ffJbNUD7MDSOj5U+PC2VaL1wEVMUk0kIoThrQpcFtWKPd3VHqQkvTSTy8XlZP
8iFP09rekVRkEv1sjzUktWBuvcWqWR/lobMUmV5Dq73qz4hvdRsRKGn/Rq7mSyIegCPrhOFfCfDP
i0s+9DvGVxJ/ZYUADu/Gg6X0h/+N6HRk70w4ZZXDU/XaAHKnM/Cu2EzHfoJ4TdA/6q88yuPViJ7/
ajCY11VAImu1QRoPF++/ZDyujWdGe0kCZ53ztbFV8u58QClKDU0qSXnPJO21pTKqgQQF6iYQhJTX
tpKoxrN3v1Fw0HD4vwmup8SHje8bCCxWsjjbatUxQYss5ZlhHkuDb6x9m4EjgnstIkE4bi3prqDY
8nP9cTe66yXgx0gMI+LyvGXHWdrXklg2NtTNKZkFubMFG8pbwD3X0PpoyYqoJT34/wmwreFuB68i
jNUWvsdr6IvgUGVGq1ScnCJkc3BwNLV9IxY/Bu0caBblsEpUoz3KyasJNIYQ7IN7YRWjbQ0XcDbo
0PkWKkhtSGZXAEKBSFAOG/RLbG8FjQfgquqzCrn334OeDCVuirHlhqU/DsnRXs2u1z9wrKmzz7ha
k1pDMxb0SDKGOMM9Sbh3oXPcBQd8wZBlggNjgce3PkmuIrfutIARgXvwxjYrpLH4t8I0Ov+Jt66B
yLJECDPP6YAJgAA1TIZNziTJqFrqYaJOApzRJic//2jEYOdL9etI597UkCDXRNiEStDBbrga54+R
9yfA+9mHTNN5b8679QOKcN9/Ji9zAgRyCEXc5SF2mOV8sHmfwh1RE8g59N56PDXDlocKwcO8lR+E
/M0bq8UhwEVrIBL/nN+H7q8l17wIT+vf6FILtk6As2V99ukXxiEaQgevMiFAj3ImHnnmE/05hVW1
W7zTb7BEgoDiy3+j0u6V9i70y1WIg9pqm0hAr5vXRNfbRxHZNoBgczC7pvQUEGgK4YjV3oOGiWi3
zBqDVRQeYre9Ec3af7DXJHSyLDHiNJM1+xnhf+tOCMRYvX5VvOE5ToTGMdQr+ZQrMtr/sHsiitfb
SSu6xyHBcIJ0sMA+Pa0PowBd/yyqOK5vz1uzlENDzuj/8+5zFBz70rAK2QvGZlkhNwCowqJ7vjhT
QWDommQ4T4WGB/N5jZrcVdvcnPgZ5492CPMVDPEhIrUWAJ9pWWRywNZMYuHDkt1TPAy6YUF2EaNZ
9pkGB28qpq7K73KvS1XMp9IjTHmTHrGSmu6Iw8KeBHiAAp6p5Onks2dZRmGqVZgfCqdrYpc/wUsl
YdpmJ9sRTxivwWOTgK5L7ALQ6tBwzflXs5OAvpqTPy4g62Iv2odmAxLOFkPOllCQjuzZ9QMITkOC
tXALvKBw68PUUAD/luKlsh2anVX0uqR6SQHVUmzkhJ6Zy55gzW233ir9OQB1aIlNv00DjUs0SSVs
abxXP4MZLqjm7HJ5P6/BThTF0cB87x6KdWSWAm0/RxghIRLqnJFVDrqy9P3gZ6vr3O6D5S97I092
UgcERA5b5laKx8ghgo2xnOLXjMZaPyxbGmDmn8VxMsOmaYuyiXOwq8CSQitoxebcrajRKIEk7/CL
R/9TchnW5RRxMdXPbmPso28rW83omUdV7ipTIHM2mUEzgPam3VNZuYhuLdgX6UtQdpE3h1MheFPX
HY1iL6xASaFAQpzOsTv4HczWNNtTEJv05DilEQK9DAbvIp2vHKzI9OghKzUtz7TGmtctR/FkN9k3
lBLrw2jmhIobJ/4lwDfSFoiGAjIu9ph2AYPDnkYlLS5w/aRfDtGhhpM+xYGRHEmI8yYI/4dqViNa
7WJBLuJrijCetqNXorK4OMqI0I+oaaCuHKFa1SCVHUF6HzFow0uAgmak3B0SVAwz0ybtR8FldFZV
p9QBO6uAaWuJjSkBE7FUxEIYfu9iqMKTXAeiOz+Lmf/i3Yxkx/rRmQOHnftoiwPCGzfoaK1xznpI
HnB0Y/n4xfts5R7usJXQ3ViixDU3YfMvYKSzs56Oy2HVc/vr/ODh1CfiVjn7lf52ZNSr3VQWJxM+
sZ1gSRxo47HxoGUQwI3daz3lDqyGIbeKtuO2ApdFY5dSijz0dH7MkiTGx7FyhMMtWRy0BnGYgoiD
3zXXt0XnkRrmR2fK8GOwWdiRlQtt51z2YjWlfgbtmHUwjaA3n+MFCi8cxDES6DM20Oks5xlRCl5r
t+h35ceByTvl31vCQaRHI4IWQnPBORc6LFJwkn2EAiCMUBDUSYqOc+d0KssMOzHlvPVnauHoIPsg
v8MC6RQjmJXEJKMngYUwC9iuU/gYSa2ttj19ivnPWiwVqM8c+HyYbn9ikX+muSHzAT3hmkF5oD+7
VF10YB9bJepLH0+1xjflvzZTKJGC4tqCcsAclCFHnxn8Bs2VrBC92W328s21eqhoUhL8bw8h+JUq
Sq7+khhyrdMMxM7WmdHd7wJgJvf5RoWehNkHiSvqUyHToHvOZl3RteoS05H0dyofn32amz9TwxcR
NN7Yt3mqlOXe9wlm1v9Zt1QZqGY+uENnEDf5aydL81Gh0OEYR3cQMqFbcjwmEhMUNLT02Zqj7Bsx
19IkrpeuUxi3QSWZAxkwz1a23CpJ6BfWXjXv9P7pr6xYDQczfrxReMjW21Z/0Y7tk7HXncYoiH0V
KNDfFZhTySiCQoOuDP9m06q7ejXOrQEbMK19ulQymut9C9gfYZAxaa2E8/Nhl2Ko4h2+W2BF1Ab4
eIpy/SgOr55ei8PAXagQDGGL9WxhbjWKKPATEYCuGVI/ShpxuHrJA4am/kPVBF1F9cr2W81bMlnc
fBP9tPUPlRHLIffWfHwdlVM7R4Ojt2zLgwk/kvv5rntw0w2jiX43t7KDG0E2cEB2FnF3DagBym0i
+eX0XUwz9selk2VLMBIsBm63EtpYVt37Ep7csG4P1OwofeF1iJAq1dw6eynaedxAVGTASAAa9g6T
jFvfoF7yk3qG8YJfmjGA8NDBIJXp9MOS10cr67xOuXvV87vYhnrstUxF9tsGOf+3RmQgvWF5TbuX
ReRt0j5nnu9ui8eZ4Q/QcbWiDI5f4XAbiB403L3HNpGPERgt75jQl4znq1Ggr+8nbk4u0nVNkqYj
fVI/Cec/rMcO4TCP3xgDKJlQQ0WsTur5whEpxGQO1ZTt9qCHZF4y/gT522z4rWLMHlc6YryIdD4R
Y0zuAMwWPYbRad/gftdqq4OT4yy+XzvPQ8iKXfoHzCIFfl71aaX7t24I3GF6NtgM17FACEZkkGzP
Rr7DelmdoS7YzhNkgMCu4tNN+OZTrYm2AZe6OgJRP/oUOyYG0ThIYM4LCjgBHwC3YUzntTyc/vJj
Ref+AfDpIXka1QUJs+wiYSCEWOahEWpDzYS3oTsy3jtYL1J6WlryXCfA1/8iayG3W4spRz1Dhdb2
FFUx5k0zlMRVDU7gxk/hzP28D1oIL9iY5A8zk/86O13G088adOvLU2NlUvHFmOFBREGjlsrG5sO0
gcb0q3cMJ6HLGnCUPRznQ0BrrgNW04z5A6jCCNKvRqXVUODNiyxbvaFklVLdCzU0U7uBWNGVJRTW
tvpxLTDXBFoIGSxoVrV1Woxu70+06Oi/tqqJM75fwAdt4V1uMNUBDYs5JHoo8rVgBG185n56yyKn
m5VWExRrB/7lQrEGfFZtg0gYLWeTUsEiWqT4XWDKZskxd08BXfnDGesyPuFSDWJE9UiYsMxCxf3U
993RAVnxwzlC0egidro5HNIRmnVXhX2a09qvnbn7fbjh9hUkV6/RN38P8Wcvtczjxa8KQo8sI9Jh
za37TKbv1aWMAHgpTrQBX38Hke4wNi2TQ5/pnHf7ZwFOD0MeHiNUVJAgHXGNhmhCv7GyLLPsl1M7
tR5pL7/zfPi+4E+T8+L1LgIcvSscK4RNnBoyTaXB8mLzFbNjbB/A8D7p8eFyBPfJmr608j6qOYyK
XagDlceGrNTgjEDRWvKwd4glPa3tkVNuLyRYGAjf2rEKN7/dePMpXG5/N7AJiYEnqNSJchSrOXHT
JUddXAaNL36n8v+XPED4lWHCOyMvVIIN4zry6pASzGt6LmDdUxg1tBZxfZLKB2//P+tYelM0U+f/
pWQHfkqHbTmUDrQ72HnynqcAPM7puDoBoVUT2Y+m6ZDFZQD94kchNBqNM6wXm66TQRsL4MBvFmBT
lOgo3Y9BkpkBD15jwbPaRBbc1JRyK1OFWu9AHL8uWCHnU2VI6ugwz3COZr3GT6aprleESIownpvh
koQLYkJW1qoZypRdIZ57L84dQTj0CzqtiE3KoCMbYQYr+qxb8DT9NhhwxG2RwmIoFplY9NiMPj7E
ea9Tdg3h03WNVtmRYIyM8THPD05t3H69DQ4eMRZCso70ITZOzYy3sF84+ACBKuAvdD5RCenCCOk2
hhoOAHTKtwLYtEfypcxAZszdTXER+m1M7ErCVtfc1+ZcLqtych2LmtcT2mtVlP6IgK2SUGijIH/l
Cxff/Ntv7K6qEEDwqAlbpBNgeB7BQyyWSOvpZa+hwn5JOViZW5/eyMxtWBMY71nBQoUCh8If2/E2
RT8RtSTfdhV5dOLwmHUWJuhtqenQbt4HZlucMVwDpFmmfJW4vIGWjz2Lh/xoXJ1/9nfnuy+J1+Ot
pIOjWhKQsT5E8UJ8OyIM/l/Uh3DuRR/LrcOKicJeok9bFInTrTPOhBZ7BHuM+mvfGSK6che4llOO
wVvgpLaEz/iltYlCs1dsfdAp93+OuvItlqXv5cQ98DVDvF1qb78AR2aZTYOGzniOLu+HJi5jiBU+
kN8EpmZCnaBiv8oz0ptP7d0vj7hIyVvCDH9cppisAsuZxxvYNulvJb8lGWLKSZ0rKVLIIIpgzeiT
dNXmahGeS4mYIx/Adxhup4//r0G/1dbrbI/PyApAFgfLsFJmye14LIAJDtzONphxZIs+G/hLVHuP
WiTNJxpsihzwAtuddIer2YX11Erq0yQLizLYFWtg2aQzlMmY7C0X5fdw0Q3PUh97ZziPrRsrTPwA
nNJP7yfxarxO8bnCW4Yrj89c0ywGII2m1TE7qpCxSOFL9fgNRQQ9TNl3S5/bto/4hKunq8D+/hem
9i6u1I1wZ7YMVph0izryZucFOFYGvD+zzR6hWJqvdQHP5AIN5wZkGxV7QoRGOUBFgHj2Rj8A8I4k
dblhkgOOzQgkC6mSfoQN/Y4awJ0LGnBfAPOhJzAQiVbJIjMV2qK12MwbjEcTufnvy2042+BnNUSL
vWYS0NcEOymzRFfnLde/1Tyrh2eQOPCdeYjQCJ5qt1W2gzOJfDMo2OTpNPFhfuePFd+ZWCE3S7a2
rJIZZr13Wr6b/gYCHCx6GrE0ylqtHHtZUTYQg4b4FejuDD8TQMjQ04+Pikf8j4wApGopZNMTxXys
ROR3ZN1hbi7XnQ1ycN7PUjwxb2givIFqI4ecTxLkUc5f6Vs2DcOskRpQhoI5Hd71sWfjEOW+Wv8t
tbfh7YLluNXwzUYVFx7xjHG3q2hDz6cxqOKe7Cj2LHt8Bcn68JOw6Qcm8OHTKd1KXTcbxvOW37p4
u/LOIZ+Y7elF3ONk9cGeFQaB4VM6waeKsaPgKK9SGPWTUUEOY1D/gUK1M/USFvq9CPsV567fIDWG
NGJCOK8HTZZJdXYLKevQajiI7zxOZ84VwFkG8XPJ5C02S7+SG4gjoJhTMH4OHp6cAs1MN/lWbb3A
gjYe6LaNRtQREXDa9w3ff3bIBNRJTWqfvZ0OHYmVjUl5xqCZ9473cV+Km44a1TK0PlFoAGqiA7W3
p/n7VbGBuPG/qNShiHAvkom4kZW66TC+5J4tm2otFLSXACzP5IHuDWgavyM+13rARnK9H8TLBnuL
AR+4FcE5f6JqaEOp2FBsGr3NMQyww2/bb63ZxCPiktEz5S7R7ye9TvK+UJv4IYtNx5lEpYOWaYkw
vVha5/XZ4yjdI6bb0ow72kX3ZnUUSOGR8ngob09rOD62tXPoK2ooqIdrrxuzpqBSpHJleZxMm1UZ
1CaePfuP6nwpQKA6qbY/gY4jEhn20ctgAQbDLw4qagMN8tMfuarj+ApCZTkxAvazY/YqBfbe8p91
2VPJVU0zbZy4Fs9d3c/Mg7eHLsgcwKVgFF2wt5P57pb8V5o0yem/I2DSCgjSP4Yly0mcK5q5NDB/
74lPXEivBH7iFrMhxQtINDrRr8a/TXt/+9Bc9+imqT7F9Q8mqJ+1SLl6Rbu6lnKlSPadBsEa2ZNs
6DsqfTfapziI7LSKGkBn/A3XJ92F1MuVb3B8ZMnso1Xf60Np++an5bIF/FGS3LHu2Qs7LDT1ANIG
OM9XrbJW0GkT0xhyUvM8Ar1kNigFAuxqbZlBq18nfDuKWgEE2vpsnoLYJHglMGj4/Q107a59pZ6a
TWs3IoruFmhso4BAi+Aftr+83fYixQ0s2/pmHH00PRFfdRUAyDcLvxtMNc2hNYaJQK7A4qxbjbCQ
Vx1mLpNGB7f/FSQgzbztu4SUNwkHKo1NFTC5/cFtrXzE9eXzjWyOkI7RJlD1zJN7Pd9jPjwxN3fp
KKd4dZilg7jrBLctHYJuI4tCdYInRBheB+rwre18Tc8jWDLHtqmzlmc4ynRGmH6jOkAhnGI1KYlg
irmgd7jbBoY/D2DGrfJB+5nUo7A6Ux65sGcmb6vPBUrV44UTw8rdestDYtvDgWWvsT4ymg4JsyE3
xnWG99eQvLGXlA2LMjsoBxZRzBytsbwB0Eu5putM0LoIoP4neYHRMW3QraUQiEhwJtJaFc2tGIWP
WdoOtLuS3Bvmp0L9z2oTXY5qKimnorSIQb5FnzUmJDTeavtcoNBCo7AnM8OzIQoQHvDCKsKCRMsO
scH8dy4QUWOe//pEF+4Cb17dwZO7RBa38pIKIa3Ymiu6c9QjsAVefsJPKc1tDKI3aoF/blWmpId7
rDj1M6YKmTrVr7YaobeqX3wHo/aRXWyag4MIFS4WTbVSMMIenlipFMIWPPUkssjAd5hSqvHSk5F0
HHoROldIls24fpuHyBzzhwHPZdp5KZmarLJkfV3FFYOYUtymQ8kmBJe95BAC5iPnybX3SkLGz/PC
A8fHGtxlBnBX7ZQdz8CfkXLAD37z9pr0lxgymcrAgb1g+3YKdUpqKf0eZy2eZ/pVW7Yy8hmenEd0
DtQhZRgBSKr2uKTDWDKj+K7ZV0mjRAVFQy5Fwf9ZP31QmjIZulpZ9R5HXcwsm22iCcQstGU9hUC7
Ht9btVYYyzpONW0PA4Jz4ipef8p+NNW9328wB3PuUgOkpLloFt37nBAJznbhBP0lNEOzjEkhcoM2
4m7lQmc3KRExAPL+WqYG8J2v9JIYxx8spsNkCgyOCKVz8QxNGYs2ivRmn3TCFGU22dgu1tS5cXn3
hQNO4iWW+6TVJVxVqIPO1R+f560xN03JlGB8lMYjvPfqi4+jzcc5lA4Q2RSGQMW71WFqcNS3FLUA
//02+nyjoqF6+jmcA8nfW1nREQrUdpopVd5AKo044O8Tx1oMJYEQ4h0o/a1HLE63s1nWsLve9cOm
CMJa++U+Gxn1tC4kwShxO4VW+YyA7ViYGKPheI96YJNLbk8ps/9l+tJxhKFwVQpsFCoUjQD4OCca
pGt0e82gIbq2UzegFeilYyLt0KxuVLibMSaLtrffdY0C4HVyg6wwWa1/LIBPS/5hE3zlkkxe0NOt
SqTub2PHGBbBhNztNxagJDTrWBNNvFzxczT66HM3JcgBuDgdoJb3BbYDid0gtyhXfhx2uH5vKiiC
EMg+jtTTqaOecWWxAXvv+zNHU+cXS2dnGNuCXZaa+h18cJLwecF4Siy7XJ/IF131vPHsVAJD8MBG
VrCgRSM0lGWn4dm2Q1vX+0f0BtTwZ9AqwEjiSL8TwUK1T8bjr5RC6YEHU9tthTjVQwXOWeO1VWqH
FGVJgY825yJkPzdDTJThbyzePLPtXkoTn03T0MIccHkN7unZX3GpzAQij+cXornZcY7m1txZmPaq
+AY3U42Bl2C+d8OslXcp3kSOA5V5KyHzR/kmukBtF5+HLl5zNNoLoiPRf64V6OYZDL9ea9L0TB0V
HX+MQaW2osJXq6OnCQ3sGhDb6lZziEvtnvENwgbgi5GB5et4HZokHX6xATBMruOm00szGYv+/AMj
Pu3BI0v4suYCSNc3eRfhbz3l0jBAHpMkTEOdeh30CZOesA+lUTcI4CEXoe6hhmfaSKbufFfp5oa3
kTVC+5uLps2R7Ewx7RLBDdxlFRAnaCZplkW+v3nAFvIULNjiEIvfDzKPc8SG8FJ5WbK4OlhCywDh
J6p65E9ukMCvYsvI51Dymvvc6icovkf4/lvFTV50uGz+SMBdjDy7rs6H+qN/BWlRzXpmj02JWmry
DHxCkfyM5zWhxUS+XxA8mmj1t+4orAMpCTrlNAIN0CpFmvFXQQ+uUj65e6yPZJ9LpZCMRtOGpwEQ
nB/1MzH71uWbh9+lDQ1DW6i1W1/FTL4WioyIJdZ18LX/gTAMzC2Ov3oQMPMWi0NYa2xOvRrA0YqA
/xtOYolqbioHn4pwngHH7sjldqCaVbIwWI+CoM3jSC069QoYfubnyLjGwkCHwGzH6oPKWNXlpo0q
ugNiwQE+FSLTpZrr+iQjw9PRJPlzWXZIt9WC2Fl+L6OvFMPwt0AF+/eBImOsDLnsGFXoHXZ1fYhM
TEf5MlOhQ49nKEVN3BXyoCtQdj2jTgfmY8fC+KzNPhq+26ejKIeT4FCGi2VW4GoZfV7teO/xq8oC
jqP3c/92b+vsONYOLalumbC5DtdUUQO8BtrXAZxxJwqv5gWrEy+sIqRXDCCgwrgbLq0CkFJRGyMk
EirJqaIUqyCr2E0OSxGBIya5YrvJPCAc7erXC9PC/cXP1yqpoUdo7LoICJ5gdjLcFlWngOTtdXME
PLwZkFgHhcNB1rMHf8Em8dAbd4bn0aoidOIhBWUYnPQ7ecZ3WxMFpvf2kGoTBqQgfEn1c+AXjNr3
we9DNURIs+qrdQ6QEDxrak5YKfiuOzb/8c2yY+l3vQGnO8HiVHppIXCWiLoywANbcSX9bt5h6g2r
UhPjuM6MKGZeZcWV0I6YWDPtX6WoH0QzraHzz3GWDXL+9Zt5NiDMdF82UG/oNeJBq2tjqvww+y4r
Y58vmSzVPfaCyFpufYiDtRJX06MnLPWa2xftabk7BvqWyiezTUbXjd7NlE3fx7lGU9iQj2Egq4BH
y26ODKzke5V9U9pNIug9TVpZpMuGc9GJDrbrSo2hM07x2ce6cLd0I1igdTFy/C8epYtdEjWF1LHF
2ViXNRb6BziJzzlRz4VGs88e2noxNmyZIUQq/FCwk1xluYO2Ou/SpvNp90rU6r9TfnT3j6Y8VP76
g1TCV8AXSn85NvRYZ89fnNWwAiuAzC0b0hKTQf5l1radVv/Ok4E34Vfva7auJ01V7jQADo6piNGE
nl2xMgsQJCYRkCZllIugKyf9GWi2Cxxh4yy0UquNweFXVX8P/21YQNi4qeXaZr+CuSg0Ra0gV7dZ
DK2JSMFcdyOhvUiRkohcklqvykxWNm40ZEzdqLV2gbb6RTY76/lRYL6XZimyL/uIKoAKoHrAIE5J
8wYikcEkhIWc3q3SMzotmqHLlIckeqUFPDjxeQq5gpYzoKHUR6EIzcRV5QkSLgwu5aP6gh5FZxGa
1yZfBokYh8z6Yt2aH9NFOb6p6E8rNYU9E2NJdb1HQVULXsMiR8zXR9drZS8I9Dr6O+vrmBqOTAeB
c/4bHRr/rfyL5LNAjScuiFUQuyN1Q3FXTNV5hf5kcspBLkACcKk5PMNiDBDb2cwrhAqZfB4nuNJF
UFjeZok6MOcQEjiGkzyKYEQwJZ/XcdEw+LwiBh3JeMWWjvNIlBEnCOFaMYJzEK4MV/iObyYBPh8P
cv9cgIhdzRWHmBIsks6RzzLU4FY85dHjy9+qGjSfMglFM89masrljpFwMUTm30liC5uU23ilaThh
QERMS+VgDpelCOugeN0r226TnP7nXxC2zWv9iYxxeoXwnXIQND2f5M55OhVj6Sb4tFPs0GkweHDO
W1REo+0Iauyxg+xelf/WMO6gfFht0w3RyEqpxp4eWubOsFTmOJSZr8LiX47dToyIEo/eMlBUns+9
tSn++0KeZeZ+9Y92lLtIvr8ZUlVNqAxhvCm/kBw236RyZp+ZCX6KNREZqqoCu/qUNpsiGr3nXGFP
Y//2fDFIlDNTIeed/0XoyLPUTvS/7EuXKqJU9jOJoHSS4KEFpaPdDjBr2cm6fPTgl9OjydkCL9Tc
M5x9zPpTJ3g6srRSv/WkZNPXlLzTkfkgYgPcYurWOuogjnZdCkGmvpdEHqODINuz9CwMuPk1zIyU
Nnf/woxR80TuUfVH1PkKn8wn9u7Gkc7hOX9iVn+2Zv33dhNutxqgkBWRpmCTqbhUJ770+MJwUTHz
CxX4ahiWNwjWIJTf2kNUxA1HHgrWXM8lDX3ybr3DuIsXCeheBdQsjz9ND3a+d3fVwlcejVuAEp8q
jFUyptNAYGif7LKUVZ4fmrlldQspqyPctHY7P8a8zRHbL0ATvvY773iZrszkCokBdgTr4phLUtmJ
q3c3Ee25NAY/pHSwlcGHXTPafV8M5zNjrnoqS8CHADz7ybUgStUfY3UmsZ9/u9Hij6UKK8F17V6b
vioMaeM+XbsbYtEqxpTyR3aeS6WiSlMPq+FJEAeUTXYybcjke8+u9etwijPzUKrbVIPjcbF6Bpp5
oz00VbeoGEpWrETXgXn9r8WBiTNNAabOyr3AAlFJdmpfrUdegE9a7NGgSuM5rGLNUUK4sgxRDF0j
tNu3EyryQFw8ZJiAkkXFwoNNhdBDxJawW5MtVdnmAq9nWFE/Rmm7U9KTPTOy6m4FNed+hwz6rzP8
Su5t7iv0oT++qwDhaP0e9kNsrxid6EljaIyE0jGRge8SvNHQ1d1/r+yceH6QnZ3/meEKo7F7lQXN
VUqcNIObnq0VYksb+SDtOg049lGb6Qzev1gwdP0fl7HO27/bn3uvFkJjEkuW0VBuSVdCdFqlMGHO
QvaVTYFnL+w8cGaY0DLK/Tt3Q0lrVW84POPq2+VFWamS0biaGcxRPDVS9KVqfg0X0KED+og959Qu
ytJEH+CkObvAHIj0RMK9aT8AufZ317fHWh8PsryTUiNQGKTq2Gqr66d7Kzy/bQlVm8WeFxYqgXIg
6F1ts5xi0HbP7uuXTDwl4TIIYFJQTBFOENFgCp70pXJdptTsqEAznETl/yniUDSEz0q742lDd/5x
HnIYp+swW7ptYfkG3KNay2u7oD/oNWe8NEv9KlLT3hFg7t2XInJb6B/i+/qHvVUpTnxwgtwzSiYG
cLWZFfnHoW0uE6rQJUsFk1E4ImYiaDu3L2SJrfCfYTTtq7FJplWtyDTGdoxmBUPmN63t3qUX2Xw6
E1wpQkyxLnY4PaJTuTE8Ve5La7VRRnJpqd97KmONi0/r5L7BePwflEGDbxzss0f3c9pdMmrT7LVg
Dl8JZ/JHD2+p/qRG83+m9gExTa2VeElsfPWZMMpZ8rsXQtXxrJ2pNsCQQ6UgB/hYlil0fSF9MXBa
UrthVG0Vdk2ogKN7AcFAOQjoKMt23r06ysm5RJd1lwX8wG76ePP3Ync7c8BJP6gyxalUB3mVpjui
/GxRMzEVYcifOCmX6uUXNTfk3jCjO6Eg/1S2Lkc3/dpNv/wJWtcpsiNM670ZJKNeO6EW08d8jjC6
ZdkAndgix5ZAMvGVtuDl0c6j3dlaiwdaf+jArRj/apoOlRKSzhvTYsqtiDqzNe4OvyeXgRsJZTN7
sVaPyQv1yVYguxSVC1oCxpp4f6pcaix7hyU3D6Lk3pI1/RHzLgzUSJfMsPYLE7vGJMR40JPyy8jr
TJZ+JN7avR0NaEVhrFoXVmjzRfYoOLQt9/i6IotuKNKCFnaFBgeV1Rb751gGCPzSuu9fhRr3eDaJ
xwAIwDuYJsvWJmRppf8mPP11b6ig7fUTa+KiaZncxbxgdaVJV8L94f//Ul3XdKMdSLm2Ctpi8phZ
VSr9h8jWiMfD6YffRMtiutD93tmTUWLfP7xb0SD4eaJVYwPu1mpP6dlMkBpK//u6rsDyOYDPYqLN
XziuuU56fq9gHIQW8GHvlhmqmd7/v6Pb68TdwfeAYE/xiJRcgZ6n7iO8Tk/76okDP0k3G8o5ii9X
iUUD3jx0CNt5qxDLv/RgkSQ4gCJLhC04pGQThoQ3tffmeleV8go53OlfsVFi/lXBxtg1dJNEW1/i
f6rgzW/0AMG3a/n6aj/EGsmya4xjT/BsmRN415lM5BudMcbOG3pbHK0bDyPnxhCHWdS60TktJWp0
+/l0G30jXeghkCp7FRFjtPyEBYKbZcNuqSS7Ujlj9J3eZI5GTkvQuNz3ffHyWaTiZEr06gYnJ5Gk
DvSuF/XmLGF/Irl5LrQDYMQ+4aoxs4gCGbBNSgX0puNFSVU/sH0dxfcw404zqGFlJhJq8/oQlfwi
MTEIdQPNnXNK14uo+HxZZ3JQOtjsiSwL0RlDuVg3rxYh1+Jkrd/NcT+KQwb+bcCm9j+dfz3oR2c3
y0drlKOGX2/+MOFOAmizsrDMKhB7LNYoZlxhsly1OGDTsua3HsZxSuVYBeEi03rHjq8Ihl5jlK4S
e5JJEhPhTjpTE1+lcCCS2sBnMZhEvIpPqqHZ+ftdXMpYwB4maY2Qj6Mdq1fXpFG7vmdONClQP826
aBEsONYDsspmuSrUHkk0SV6+QgOV0h/taI6vlkxz0YfFSnUs9bdUHJL2uM4eb2z9myaYXhsozHyj
CmLuNrXZv+8dkw1MtMZMWwandlZZKjP5pzulGllGWGO8//f4uytHzsM7iNV6bhjd+Di8JOs4LSfQ
ywCsdVY/OEzjESH51Hwd5iGCrGN/ZqfKssybTH9yEwYOeVq+qYFGaammuvzdGReTggDQ9Gnv+SFu
kt8QYHFqdpuhHI+IZwExWxl50zNtDW27EDwmV2tLlCs7sqQQxFbXAJjm7csglfp9IJdWlCBBP50/
ndNEkoqZBQLvWxZqvAHQ/FBuqddH5TC/ooslCXx0uCAugrfjo/ZFG41kmaAyYVSECB9LqDGUvTJI
haZf7pvLYljL/buKqooVHKnEBkdyJI0/gIieuapM+6dxa85yg17T28afbTZOXZFhtGUNKYUVYlMT
weLIO9zfq239a/1kwcCKc4ym8qz7TtpvaL9sd35qh2zdUaR3wZiF/9tStmi2lYbHWe4ykr+gHRQy
suE5AFNw5tIxi1cryxAZ5zZ7sddjmIxg+FfTnwO9WsJ/OyzBnQnHI00+hLIxAAfro4cjn8FcaDNw
sFRhNns3o6bpl4QFL4A6Rw/Aj62Sx+IN6dW0k5P3A3j91q5RDFCxRSL18elsl3PCaWCXRbz1ta/h
Xe7jdeo6H8G5KxDh2UOhrl+DcHMq1NNoKJVnWhPfa4HDqaQhbHyT64tbHbJVGefQdFi24y6UptTZ
CDLbOhhZEHJa+Z4aYW+HRPm8oQcFurQ2NiVZtO8P7BuFZx30WiV8yQr1T9evUUi6ta3BjkKZQHt3
YGnXlXv+vLZkcfmlZW/QBgsKq2+fFymkY7hjoyoE6g4y+z9bBQzw++zkkjxapS2IcmKV75g+cj+1
4H1/mrngePgGtq1+rSy+G62FNyLl4CZ0CdY3gYqitVDPbHyLiYX5YeNrkK3h4Mz0psQqHoLLRB1t
qkwt6pwJJ6PDRjc2Je26XOjeWzajZsQtBedJNnRY4NsvQdKW5JpWbIOuZoTzHXovCgS41i6zHZD2
SCCXlyEQe/3GfKwi+3mQd6qXRaKYn0MH7Ur3sH3hBV2nSJHpaabRSBPAqLWDvlWt6FnByitrtGdf
fwHxydP4sBfSDxp+TBbdZqexpGeMn4NRmR1S+Wwf1Kp1w5i3O7JEaGPspm6zhWK9hW6ShKOSPHD2
ooC6rMtO4EnzOnkxwgwhGIYlPZ6cbcv73oyypu0SSl7n/t5dUcMVSfyBd4JeVALMfNnysYZc4Yy8
GYeSdGUevc32+cdWi83CuS30POaxgSWU+jt36af3udsAvtkFhPK6VQkR1PkAXAmUAbh8r27wkVpC
Bmjmod+9MM9TfNnV9QWhajJMFcVjdSTJVbw/+f2/bWClQmHMtxC4FXJHaEd+q4F26PqRr9g6IuMY
5+u0aq2008t2BWZ21kkefsZb80yCdsnvnaTGjy48zO5ZhIKL8pZPFdY8xR4hFSZEpkABBjB8ToCm
d01x9s+BJBVf5co/C93XsFsanoYCdpgulcTgtahN4iUela2TSl1Kn+/WhORv9rYTjSgT3GExLK6x
Sgx876f1z3DCaRBTE/4pI6Qj/KOlE4ECNnKBSFaA6jpsn4OEtileYw6rS9V3PwwU8/y6p0MU6ABQ
hPnGCj5vIq69AJ8perSong7M4E7x9EcC1WBX+lBFeW1noJFgruUg0+i18MZHafYvIuT+NrqnEwb2
tq2HOgUwZ2m/Rw5NYVoTRwFSl5Y9eOCYE6YyQ713nNdIxfqZKkeQO8Naw3W0AZLFKDUfsDNvh342
N4B7bS3opFQShUTBw60ePex9/dKg25s39Do0M7ErmKA6St1atrRtQnm5Y4V1mBxZWP+LeqXQ0zTU
Rr6UAvyYxk0YMjFY0rtD/YdiaAm0v/NEm7JNT9FH7OQG9c1x5DfoPCBTo6kzOOlXe4NN7rrk2oOi
UQhoPy8ExvOja76K9o8EUT29ba9VHMg+uNGZBG5fKeRYk3pnw6C/4ywDMHkqEf3mMTLWysNiNSXM
5gmNzj6xoPxJXMBYlq2zjfcgf/IsjezBjLZaxybnA/LezCe3k/AWywRQPWQfDyS4nPybcBR3dqZy
rChKRHGW2qku+0I2QvCP7SHg7ICqORwcVLm/yJeOf547/TJ0pR/71ggUg5fgNhUBmM8Wfv4vSMfa
ccYW5vr6SruDDMTSjH5VIWBF71T8LODcWWqYUkms6dNsqrWzVXny4/16AsQfE9u424b6rINMIYB5
dA6PfWw4WEcv8hme57zOcC/A4ScSN2V1sqe4Pi/SfkBtYZF2DuI1bBrkuHpfwE764lwcoASkb9bj
1hnj8iETodc4ia5QtyHRq03KkB4mWImFFE8LgwZyeAKkEAzqjRUyUcML8dDj6lXMH1qu56JTmKKw
11Oh0aznhm0Mb/Aguo4UPokGFB4NTfxJ/WSLykuoLMsKO+kn5RToWB0WLLIJgpMOwYK+Tv5vKTjw
RJWVMjPI5uOt4VUAP+nDhcXr0HG0xc4dTKwMV9ktfHxsnP6xRvv1kBY3L3wF/KbDKWUUihLN0han
LXb2fF7khed2i+0Kq4XM0EVH2zc6K8UphTsZS3zuTIPfdnoNcqzxH+GVMqNtnNtBx66iFKUFP3FI
qWmOpgiCYLLuCaXVlNNj/m0kPXUGt41X2MJueB82Bc1ANgZYpe07hRdCq+ltAlMebfzgo8RVSCRf
W2aXyhLP50Jnpv8gCWK61i8Ve3mtKfyrhsXnMD7u1vFwvja/9OJqTDMXzTFYRFvtBE249E4AUXwN
V5Ha6iYusXTJdW4sWFZsmJrmLxIFh0LXVBkiKqg7jgGMgWtSw5XXdTJ+Bqq9hebSsjNnvczVGou6
HAKM3HY2wlOX8KxfYyXgzIwjt24Dl1uSZoZ/ISCGqGjJPgL8ojpDrMjpPcvfHcIlk3DZf8X0SY3r
W0VLBw/SLvJdQPgMHd36FTUKxTC27dX+KhUGMKRl+J8Yg+NC2Vkqn/uvxGDZ03poqeTDYl78ejGZ
QNnKVzBXacrMoYt/N0TDMVOtaSRWZD/tzbW201sosag4hW4Asn+RgrJb82LTg25L4om7UlsW9aXp
wfbrIHuwzQhA99ZyqVkGpdz+5zdqV/c9ak9RF26wRrb6njUEJ7D/n8UGBfO2f15VZYfNdGI3m8W/
I9TrVm+SDzhYCB8Ok0rkfdFZTTBS8J7IRJODN1tCFRqBuj5nU4PFJGcY5FsOjwu1DauEWYEzILw1
UQ9uMXwZqGU/ke1Of0+f9kflIAZGZ+78eXMMbIhajwfidOky2C7JS4wW6LkZsa9tl2fmWG90w0Us
fdKeERmV8MIpRa/IPld6DfWrmUHF4FvtrhQdcoojaMP3cs/9V7Yw6WQAbxfFuweXh5VrMNJRNyk0
MgiLswHIyBi7WvoUH3e93u8A5j3POSWKCN4tJ8gIjrDty9StgvOvnwQnMTDe50qHk6fHL/aoYlZ8
Gj4GVqrqmHdMQlr20ayI6ji8vn1mgIpnNvgOfAu+KH+vzS8r7En6loIBHodWvyiIP/S+KKien3kQ
pt6j9avnsZ61+f8HjFx2JdX5ZsANJpJHnmsMoCzWh5vSknc+J2x+Bvni4yxiF4ULd6MYpS6EZXdi
MFXUNIor3VaagNq0zQBoyYjkM1WRtRQw3Qwnx16+hcHJs0SvLxMMjtGDTc7uHkLjrC3sqHs/c9S/
eDNzWub5wknNmAMReCGM+YdMlBV+X0b4E7GetkeBuQyMUYTISGvBC181wmfgl2hIcl/lj0xHRzq3
8JO2nxISV/gNL2rQGrdyzfgA1FKdOSTQOOzPn0EvNlgvl/bDK3/X7WHPgHrHU2/QUOp1qDNmRDtx
0DSKqVwdZ4+iSjHCZ76Lsap4I8gybGXzU1+vMac2vadLDa4dlnHMpvuSjnDqvfN+NH7G2akXSWKB
zo6Wogbl2rcCuUIppznu8mUJht3vUZssBQczes6AYQTyFFPCQ1U42xqlClax5RcEo3V7Ck2kvETD
xR4N0SH1sforHOTLgVM6u0rYZMyfgppVw3gG0/VC3Ksqxua/RnGJTQa9hvtH3z32/v/iPPVnPypz
zqYbSTi+H5a6gmoUV3w/GAXtIvcLwXt7wAYJOYVKhtJJM7c6g92n9XrTKX5NS/iIVnkTEzkz6XV9
VEqB3wbeRtv9d5RJ7NruvVSmYIaxZS5vJjYp+57+NvJ47hQ/zYcQNCJiTSfO0faVJp20pPTrbc28
tYtylc/3AKJ5XUFO10M3QZalvhhnZPownrDlio9/KEh7VYqBcfEgjaUpxVEu2ECcnZMdTw83Slpm
5FVHBllWZyS7XLsLuTZZ+EwDdwpy6ESIMMVCGMl/wn025hJAPL7t4rQ/nU78bvuOSsCvCTNE0Edo
am4XpuPoV4whU8FuSpQxOy3CSvqKYsCqjtUjRo2bJkvdm6E2vlK2gA2fs8zeVUh60jLmFMyYm8eo
RmoY9Jv9XAH2LwD2LvHoZdR58IwJNmS1/hTKzqtvI311dwH99+i2o3voRT0OJSNL1FdAiYA5Q+sk
Fqx35FTVPLzu7DW830CFbFNOnhiPMKC1oeQEShHm9ys0f1GMufoec7re5I41Vm4SlVMBJ+JARS8G
G+WfoZl3svaXgITj+ydpF+bs84KANUkiDjVY2vuRi/V+p4739qbtq6ExABBOruJtY068oBZMRRph
kz3kmZn2E1o6xvEuG44cCrYdxYnhfjOGgAyExtFI105uWU3KbVAJeCc/ytz+afVmL8CEsDedqziV
rRnQF2QNLTU2T5LWsPePqRh7bNm0GZHaia4YbukmZ1+1AhKauK+rUMkIyZsX9221jkkxmLh1qpEB
M/YRGJ+YHnxZstT1i5s1P4V6KIL9rHDUk1eKiI3FZ7fIYT0Tgq8zSUAoRwBN2tjJdZ+I9gBDGK3e
P8aT/oRR9rYK8AoL6jfVc1uElpzv1BEW4cTAPWJO8V4xKYc2PriT0pxbU12pKQoFrDimSU2NKVh+
angWIsawPIX/8XttA334DgybCyjgeXbTbF2yN7mJGdOw4SFsXXvW2dxk5GmIbCsssSGWskjQYTZW
5QiS65nqX8bDf5DUn6nJ22sq+wptPRVWDSCQdB2Ji+JBsyiab1ytINADDrr5UGT7VCu+w6VjrwY0
X9BQ4ujMWI3LfBPKPpkbrMY30NhOmpjCUVHeXiu9be3WZ/T9uSJUAVatnCIF6d1N0D8afyIsoUGW
beddjBujyhflDtPxVFdxbmrmy5qiNbO3JyELIbmSBZnk+5BOlLhjBniLQkWnKhrNT3d/JAYiOiCW
tMgY8wddU3crGeco2JKA++zFC1ZVH1WSPlbCmEtfrwaG4nUuaGpagPiUI0u0ArOqvJziwrLVZMaU
HCQ1MkGjZjjmPdW7JLgVY+JJSIWdSDcdqFw9PqNnvj6ZoMN+mq6LPR7c4lAkmECAyQvVDi1LjNw4
+EYIGIUjfp7LOd42g3H5+llVnf2rHF8StH0CZzXwCo6KhcVq/GVTQrkf+yCtLYYOyWQrXiu6FGoX
B4s9kZtw8dYKUgwtkRTVtZSNQxasuhr1Mz/wxOe9tTLQoln1AZoVD1h9UPdAtA30zrASizM+JG9f
1fLrqq144n/1pccLbmEk8/V4URH+ElPKPnPDBVo9msu+WwTJbCoJ1pwbOAtSc34LxGp3vE2GFuk6
sm3gvvfwwxvErYC5D20HXsj6IgqIEkz8hY3DBgrMICLe80tUrdhxfzI23UjwE5hXYGZjO4Y5ey3z
qmrlBPJZE1rCC/Sr9+XBQ3oer1gBbZfe6e3JBxpPBuE/83QGn27KVQpFS9cWFTMcbhYSjirBN7gh
/dIrSkRdnWnEyyQHPXu+nGmDZQtIfa7lNfYrYIGS3nRpolkWAsKOa7ZUDwDWA4XVBgMf3KNuJuwm
hWHdtymDUj+TKv1vqgW53KOU99rTZfUq4XgNY7p1M/cMM7UzF05NMarYZYKQpnSMOrD0sZaF3PRM
yOwLz8ukABbP93owcZDQniSMmCpTrpLk0z5gy5W0kCKRVdE3JuunWK89HJlvwdncJp+Y739nTKvG
QIkCh5Qn9AfHtknCAJw96H0ggGZk2i/gOMmCrBA8wwwgL5Wm0QOXF7upWo32XCvTe+Gf4qGuk3o/
iwqP+f0lBrA0woOclvh1s3qPv05cgrZdlyk4pYJCNK7Com9D/S+D12qsUoUwEXlPCIr/Ttq0E4tR
C4B00YQdN4cgUQIpWPYc7CVbnUZkT9ONF9W7w4pVeEfnim+kndmUqCrIt1EICnvijoiQaKslhH9m
/Yly6U/8M6w2kR7IIiEZOCizW6Y+rLO6ByBbD0Q6OsQgrMbbdk8+tgJ/Jl6kR+NtFXIytHQWV9if
F9O6489fBVhOAGxEEzVOny+q/+BPq384qlQ3zORUKgVhwfFVMbEEb6cMhYSm/TblY9/OL+kyp3Hw
llN6/DqVPk9YZ1D627vKPY4y+P5yxZbKNLYuVGJyprxXNEVNV3YbYFPeCIz1BkLrU2JtD0FL4NYi
KMZviVHgxisEjK1RpnFGQRwR5rKz8f6aN5X2ECRJLpoeDFAf+eivYyoh4g9Gcxm6GqWH46mgPyQc
A42cW9RLQD8FQXgolOF+4cn3e2Pbs+cmIoTFAkyv1TmMn1zEPu+p5tbZGC9h1/lBtdK5WMC1fiLY
udDvHOXzN/wxpTt2DfjFL0SP7esTavKpvAfrWJ575wfXH2BLy/Y9Q8qqJA88o43HA0YsBJBIujFm
4cx3O7wteOWTX1kift9D3QbKEquZ1qYnixQqKRhz5sd7wXW4BS1XCazTAYsnpKXqZvXnUtjRtl8d
nKRPEUP5evwewlEcqZmxwJv/vvK7tj2osnRzBJpWXray9q75pin1WtB3lIUOcrZ0euJyRPJVyEkY
HN/Dd+tbj6ySNObWeHr4SIh1GQPocn7UPB8/ib3ETWyFNZWqH8gitSX7yiMSlhR0v268Lg4XFWlt
uOAxNAMjZaCan4BIMGZCXVjdeW3D9/j9bIUhn1kSSpK2aUX5IAy8cC7qlOpRYcUnEqau0BJvv53J
qQLz6PumTyhsfBSeRt4yMKq5Khf/4c4CX9Sy3/M+b/GlsvW/mBnecsrXzkbc8+We8/pE2qWNlsB4
CVAboDPdiWV2JWADj1Ygjw0+AgMoUtYAmvhg5W3OI9Ol4tnaSXwANQ8OnnBfbQKvtMBWufMqrUnN
wGnTiNm69hw2mHq3TcuWa8bqYdQxDr4ekMhrcQK59+WhKzuFXfGCd1RfZaBpmGlCWU0zuAqnl0VT
/LF+dVIJpp6nj/7KCz0lpKknx7zh4Ya4XBk58K3homtfPlLny2loy38Z1yTWT5m+mBHIfEL/r/Ws
zoZbrXhabNW0lECCxinYH3KKvci7gTBW4kCqNkd6rqvOzdFnTlmRMBTO8kT2LnH+gb9FoIc23pdz
Lm6jjOhUE4Jif9B3YWaVWHmZBFxuD/7mLFTUPqDb6MlKBio72bfFUvLQ9LIO0MztXKajuOoVHP+V
hjmAlmrVImuDn2C7g/hPEv4pMROGW3XGn9LDZ8YcZgwR7gZFVYqHyTc6tx7QnySoNTzr76R2ZYr4
G4qPGbhR8QeL9oK4yGrt4kPtVbgRHdBAPAPQXfmkpAScM72s4EkfpQ0VtqZK0NqMjq6DuRXBLjl6
2tjltoSAc7h2JfgJjDxsGpIBOPajtDFiyrdhT0VJ8HwHon4/CX+2+y00M9CeZX2kNNBdupAB1Dk4
G7SLT434alnAgy3legOZLV+WUmJ9+n6/vx0gCssGmH4ixPalj3oxB1+R2+9sUSLx49u9fXdgWpR+
HvclmVnjFtedWKCyKlrmVU+W2oG0WPSC2iSdOOVs2OCBgkKiAPUUyhHnA9pGtkRI613exTIS39SD
zC/gv3oiq1a3XrA3lfFG2Y4fLjjWmetu1tJEurkf7eNknRT/7YWhaC09ZzeBOZD8BONse8Wrjk9N
3aTN88pidHyzV1IiHdZHweQn0/YSwYxxramWG+Cy0KSn957dBFKAQDHjrgmFzdwq2FfHLKWOFmPF
ZZzrcJPAAb4bX01kXUPrLdfy5jlugHNnl0gjSX4bom+YS1AB5yLL62/7dT/KNtHJqGFw2dR2aBpZ
he4sc82DwRIqHbxo3j6OB4aZu9U2/fn+4nPNVeHix2g0/G2sHI/dN75M/x9ZTfdSQprPZN70V8PG
LHtT78cvM6F1QHmMsrd8EXY9pmRl8XmAYrqA1ryISdFg9RWSMiJgfJDooQRBBjd3duxPU/GPDc0i
It1641r5stuxf/zuunY7kO3s66kLueJLMyppspljrwn7nP7rps/1ntOVuUghx/q4SpYOZGWSeNm3
AyDmzAibR4VAZjmlwXDDXmvUzC1AZ/rK4+sPYahnPvq84H/3NZJMcczf/ghKmjtAofhslBcrCmGE
K4rqcBPVc3gj7ynS5zPO2HHYE21QEBbpxjh69fVQOS2uly6//DhL2ZOXrJ9Bt9Qpj9c2nUKjUZej
0ALdO11sKr9+JwJGNZatD4ghnVvpWxpwXtymiv5+Wee91mnSqO4vqqzMryC7I4fffCM+8iKbP6am
SGQexJf3XUu6+8oRDgEZtFENCiu7EmxYH8OzBy7HcSU/4WPj8a4g4+WYjARsMza88iuU2MJlNUdB
2UE1SXeVKKv3OmftR/c/5UtYCl5IVeMuaPmNmA8fEx6lGMUGlipvmiDCS22DglnYGR8p8L95NdxO
hxOTasAbZG/JApqRkJI3FaPNXeX5RQGKk8vDsI5eYlq4wOSi2Y3e8QfT+uXQGtbWcIDOHsbGouBf
eyCor7vlqf/VGS5R3ZHz9NKs9mj45KuBPAfk30aro63EYgv7SFviXFiOuSLdKsMrWUAtKQ2xbuD2
Dgfe/pHVhY509Kb+M5JsCVz3x+Y+gxHgVz5LCEdqwZ781GmcsIki7wgUcE0Un5yj24lzGvhObVK+
6WoI9xhFB4DR13T0sjGeTisQK95arcb+DGNPOePcU2aBu2bCxz8oz5MDzv6cPAHVtOmwlBYqFdCf
DjpaddGpheb04kPNJs20Z8883dy2hV5YlJdswMTXW7R4OKvrKU2D1RcUsc7SO9ogfoNUyGbWBsYW
NeAAwT1ndTt78ahBSHzSMbhi0ev/kV3IpxN4N8k95mUT/iyG2WEolA1SDwePN9ep8V50VNIY0D7v
ynqKDxOiVhN8U5IomIyQ3fGETgs5/8VLcLClSkOZOEkadVQOhFPj/692SpynxKPn9bUrqNzdQxiI
qdUKjb/2uoK1hkSCxEGyho2hkB5B9uEM/PPhOaaPQvurknPeMccbTdas8DDd5x0WVCc5lIPcDhse
O0dteeTvtdAFrzFgPSuVRIoDhzg5MiKQNW4SmL3F65raXQDCFWVVIABrn8ogAVJyuu2JX3L1nbGa
7qqSj8qzGjzr2OFqet+Y3TURMRcbQx/jGQMFfbAc0V7Tkx/yFP62C3p8zgkhjKXjMC5FMM/P86mh
Wz2sud0Eqi05Pz5btsiHzXitCv3Z0GI8kbv+HzBB93TfpVfV9AB5XcnUYcnfy3mH5l7KsocEB8LG
kjT/HHK+NAxi1tjDRZ4MIStOZr62/n6kWRTC83OzFF/ONrZkjqRVtPqu2EdU1avTBZuL1O1xKZl9
Osc8+Rz17wLSF6Azz49ycL8w+iUDlMiBFrctpyPLrSidxsdvOf+OXKgCuDoAkv8PgagSnX2EjmU0
jOCGVm+7BDctaBuq+FaJLtWevi7LwdT8GJqGxCqs7xT3YIvmrsCHbABTf465ZzIWpSVC+UH70pDg
K2OgItaSS+GXF6IB4WpenRhqwTLgeQBUL0Kyq7pJeTIFMdu+MR1ereTkseEw2+K7Zd2I83uGEREI
a3hr+D8aJCu4mUw9pwTvyO8izp0sbRj5chNJx0cX3Rc77vXlDtaHAwshNbqU8jexqmhtwl9wcY4f
UswU6F+h3+H/MUtNtvbx3W83MYPcmOyCSZ6fl0pIg17LfM+oFOgHJcmdzB9jPY+evIYcNnGgYv/z
3rvrf5GBmDYNFzCgC6jUs8J6K6f4qz/9bPydv2oRKwJuQiekvuXsUda4IeLDa0KcIJNA81BVvExl
Z+OYB8ZorD4SczttVc8ea0WolpoSrX819JBoot8RN0yNDRFxja7DL9mMjcKDSvAqNzt6Ocwq6Mg6
BI30oZngDWR6p9LljKJ7W2FDyFHMtMlO4j17doGeCTCidV1YVSknssnZc2L1MZ9sIpZZluBINVDd
gh6suy1fbUAVY7CY+J9KlwYl/P2PVQnkdXS/bvagURtrwiHpTULCIO4TAh9O7VH1phajmE2Qz6O2
QmD2VDBWKSXmmx5aGU2h9ZjpawkWjfXwZys+6JuJ9wvThfZBPjmP20k1kqjLTwtCWNYXgbSoYGEO
iWbdY3UcR5KXG+hiwT/k0p+Nrew7VQxp06lAbogNSAGjU+gCqQAEWcVRCJmstEk5gJ0bZE/srkwJ
nX0fpdrF/X/dhh3MNDFPK0kmfHpUDkaBbb46a+Iw7XSdayvMVRxzLJ3WIcm0e/LMGrtiZ8w2Oquo
p9HypjRiIamdIWb6UyJUxOMcWOoPWmEEk+cRQ5crS2GMSOp0SO70PCSp32Sn5pG0adukXkt8zlDp
Ic+Xuz955pJ32l1Y7EmJsBg0z2ZyBEdQG4VDhEfJZoHOLEAI5Ilz9fW0uAZLonCjqkXhgrM8vzSG
s0FI7CAYx3jt/Q4jIOTEsPXpdNvZ8zx+vutUdHkxXmBR6HxY5u+/Vn0TARxEw1sCUTQJAOx+BRzn
DbJTKFt1ARiqolXfAhw60Nf1szbtQg0wk3GBu5QU2rZXHuPSFfuIZmtOb0wNDKORy++4eXdlVV12
V1TnEqtwW+Y/TmFJddltNaRiDPGoDe+6Svux16PK0Yko5x8IRK+VJMRL83xx/+oizkEEZpmu2Apk
TlTAdo6Y9I2LYpKVC0WOWqkjhOv1A+5+v3zW7Ak9jdBCwacHphe9L+JDDB2rhpxykFMylW4b7ZPB
ysPYHA9Hi94RCnIsdKVVB/6wvSuZzWlqF9yUlsAe6mUrHuoXfASDGJWc75H6CfRpEIHDVNzT05bf
bnH5oyd2rytg8DTaO/wF+blltAPWA+hAsJQWQ5Ge9YOdVYq2TQp1zgowbF4Dw7RXbhSRreFCMNL1
kXz8r9YBgdMPVYPPDdIqGSfFVR35Ok2OY/QFgtys26bYb34zErXWjRsLcHrmSK2m+CbEA0wKlAcv
ajSnFdT99GTVFISeTUxAU7vrBGJTTsUtT9aMJqalAl/Bz24nf9HfxZ7HJfo6B8WqguO4S202Sobu
qr9cJq0i4FFRohH5Fi7QsAYewHggNc2behGXvG6BpAIXOTGvgsIjsS+jDg/WSbjP1TQXff7T8W5k
P2GxSTXyqnAgarmTOIMe+j+r1bTno9qfp6QSWj41XGtDljFp3WBbIcoNMVtvR/0n/+/OmuRKZ5+g
k7Ljc3xcxTjfjhIgw4I1YD3MYjeUL2tcmqPQC+z3c4lmPEL1JYxQGnBaYz1OrdDOptZxoigmvkeq
f7YbmZAIsbfrJPWt3UDVNNw7Qf6c1FtA3AyE+PBQB178/e8N8VtBtEDYT6JFD5XeEd4qfwuMgeJS
D1eS58l/BqvhxOhdD2mAm+YvxeyvkifkBb2SDNE5+bphB8M8pjgoATGWQGGcGfALQUNmgr5lP7rP
wbHAefGh2I+VPHjZJ33y+5/8mQMsQ9EsNLo+dedzc9gCs4GvlbZt0Krv4PyHHXAUorYdEyGwM+Xo
vmFL6cUFvhowIQqxqm1yVXphw3qB4A1OKZ2GHkPRLR4td0K7UZzYXikx9i9533RS6tvokJQPZWgH
050LhmmgqjQDEx1Ho89bVgnQ3WtkekX9PWRuG8+BtXInzAL0zb7CFEnFZVQz4pmMXFLliTJ2RmLw
bPTJ8QGZef4jc0cu0/y1KHihtzHNejN8TzBoZE+rnv1Ad8jotxq7asnBsQjMEqYnX2Mbzs4YdALU
cH19/USWtRngzuVJcrhKjoccWB/S8/wVARVRpwi1sczkhqoONGOTo43z/28gZ3MfpKZrodObdeGJ
OyL7L8MQVK6C1SCae2aOVj3uJPEG91di9XPXF3u5smPjJDK5s9CqSd9XkiblTdupUr/WSSEH3PG1
X/yQ+jQbdayYveHiAjBCLoiEBg5BBbVNjzUalLw5gCLW9GxFUzBwUFKX7JJuoPYuc8OOOdliqVX5
mbn89I2997ssiFw1GcBd0VCkLgaPWvzrCwvokXJaltSwPH4NDhlPHcuuSrk5Auv5w7lh8gn4PsRo
AGxKmV3lDecmgiZEQRzptm0Xp7poyAUbAQ2/5dowZmttGRy7MSy6oskCHNVmV3Zxh8m2XMDsJ4bp
M5r05PHp2miQUH7m/PYoZjx6WlywMaZrub8xq7qMwQvqS9O6LF6t82He0Bwgcenla00jd+BKQiVA
1E0NpIQxbk4yU49neWBqT/EUdWj7TDs49WQGktXoFhuzfhKPArfe8tmFWfSJEfvX644rNUc6gfIO
e5L6b+zNh0Tbi1GIOy5U9cBEigbJV8PncDNbcMO0Qb0SyHpvYA5kCKxDjVUlTAeHriqstPf8XzQe
FPMIQMlWVtZfKwNjLc3O/xPu8R8SKKsfalC3HquvP0yn1UMcs/tdfESxsjR5GRb98lM9zZnmbIuW
ZtOJG40ltJaUansRe8xMq8Jpg6W6lteN+gTEMximuey+YhELtIcRqrC1+vnA7lNLr5ssuI09mgDm
oicMqkFZnax7sadYvsXV1J1iwZPqH1Q2oy9RAxSy5pbeH352eWl/h0JF/i/hXzPtNo/s8kjtamwt
YKqt+dbmq8BbgnqyWkjymSM0dah2eUu7lB3aJ0c4tF4jmYc9s8UbKl/Xuot/KJUDkIzc2c6sT91t
PpCAeqJELYf1eh4MGufvPTjulqpq6FDhJuFRh7haTXoKQAY1mYjB2z6H/9ISOL3uDWO9IGqb5sKo
jLKyusp5iPw9s5IwgzGveHnkbbQPk5g8L9mZRcPtDlZQJt0qodfMGh+bILK5UXfM+uljlErPlxWy
TyJmKmQQ+LhB/aWchd/X4VeKkffCexCh+CGiwT9fJl/Ss0xL7fDXtyqh+bOn++meZ3mjnsvhXnyT
8scwX7kMV85AHks6lK5hkYv7mXKcZHcH4qGs7NVUotGN31paGfTr8/K5YaobjgrSBaDvzr6WeXGH
rbt1CLsM0QxGVJGDTkqYiX0pxlZTLtC1eDcUapqxfDBQZd4y5URD++aphdaGwMURTkKb/Hy5BiHy
7XKcds7emN/VbC+BMZ+3z1n8r8pmctTL7ils9+GgFRNtsYbVQjH9reBw9n/VQw8/YzuyBBjdV0UR
28wcaaiFc13p+BPC57uyENeQSWTyZtDyWnRvZbCPBP9FJLYWjLICBHf+xXCKVsuLgWc1pGlE238n
WL99GyS6wCI0+QSlrO6lTgneSM5DfOMc37dW6qtQzbB1hIiT6W34b+scFX44kNGrmSx9+whqtB/N
QAQVWoNyw/v9Jn8jKZWIyxQYNMf2WGhvumwB+GJqfhBt6b8krgK7d2ARqktgXEUJlwfbxmvuFxWK
+KiXb14HnGdqxYKQKpim8WI0z8Q6NNzB/mqkPJFpSZ3agZhlU8BX9pNBNjB8LL8Kt2gX4GI85G6E
DymBGfoZrsNoG4dudQDNEzJSUlCk+pkndM1ccgESC+hY5IFQSHthk3+tFZPu3O7jD8W7te5CPgV4
nqinG/qlHZcjiV26b7RHzs3b5RYi/ceqagJt7JblqHl0Rj4+k+DNGRgDSyuXFXJ6GqwbKk1JVUum
7QSMONiHjd6k6EcduQ3YPGW1PKpx0xJPXWSEDSaARrOI496DXZuZ/P3aIzk2NXlPxG5NnUfamu3U
5r8XXZzG4xG0oyKUS7g3ZoYpl61yWmlbrafvKX1vanD4BmvIROwWLp85+My8QpGVvxdJH3csB1kf
BE8Iij+BlTSXT3pgQ6V4Epj28Lq6Il/bsf1/vXL2NYqaV35pDYTEti9ex25M+Tc9KIq7pMfJ/no7
w3Ebj2foJHhH0rK1ec+KV+shvNTIMmiIBECi+ov80yZTAztYvHawdOhv/dzrlRMGpInemuvb7Wj2
vRFlmjw6E/UgR6wK1cgIaqdBVIVVT91h+E4BW2m+Jn+g86/uLuNc4Kp2ik+PK5VpG0w/0NPwGblG
UQHJA4Dj4ie2ztgrk/8OssU7bTULX7/l/q2b8e2VDjsjPMeiyp3Re9c3Tean/IKRWI25mtY8eM1U
AQc8O3PCEjPQAXqgTUtrpTgqLLryW72DlTJ5YzRCRTbhKj9AOCXsP+mpynZiYrCs9PNBYr4KuEWQ
7d2ngnF5ZPZiR19e55+LQMPZnlWvKiwdar/SVV1q5v71YSmbSrY/wGxj02QGX+JpmjVlP0lXvvsP
t/VHcsWYSHZlhWkB7B5Vq29/5l40T7WHKxEH05f1s/ZLZjZaOPKGulm9KhBXiPrc6L2GRHf6/KsE
ZxOtuf16OiTmNangAfz4Y80/23o5GQF4huBa5SkwcDWhANDLTC9C0c19vyRC2cUxPKJ+4qfJG/nB
sYdmrUiqZpuK9oR8h2V53f59wkyXVr/ooMMSn158DN2/FszIprBVDc/t3W4hVRUWKXaIq2TTJjS0
Z7DWXautrag3TS6J1Rw6hs0F6jnp802yaw8d7yPhe/svEFOiQ+FC7WWQShVlxdo4wzk7afOfYnRE
MqXaiCAO/S8Tg3gWM1vOWeqKYRVgvibPQI3MBeIq+sizTPy6QQllWfpgy/MAA3ss7lXtyON2s4ey
YCFdgYVLTvZBlDvgmg34cZLqul7EeFjoBgD9P6gpnB0dMS9dAxxcnNnYNall7aulMf5K3juITfO+
K3nU0OaRjZYj5uve9tpW+oar7UJmdnNRPeMxIOZRap8zUpYnjsFilyoDmgC/Dq14oclFAy5NPsPa
k8AnDJye3nYRQPfBeOWZkn9RPZh0ljPeiiwK8NQJratO26ixc266jPE/aYDgur57v6VecgI13lZC
+lOvEKZ6+6AgiDCX6Sy1LjcS6tCvrh4EPD/4OWmGhj9NvmfZG70+czb+0yrujmyaRZ7bTNGAEs3i
Qip61Oblr2oONxpchoW6inKKuad9Pw6Mxw5iGDrjQiKDAt5VhOshhHAGJI5v/7NdOwDn0XHpLHWk
3wUm+2zUvaguwp72jNoZ6BlX/O7yx4RDLtT4SCnEMeU2/NfMZjCTiQrHAWV37rO53xMLrSko4D5L
C2twiYQXCecthSSH3JKUudSW3UBhgEXPEi4SFhNQ07djfYMzhpX/frnDhsFiRa+UPENuX/p19Mt0
zDIR0M92XQNQuJLSmnCg84r8r735c3c2AfUmQg/6QLnAPY6geEkm7+ZNOqLwN34fwuEKhgpevaaL
FvgE77JJk8g0nboU1glfyWPCadNd5/azxshuYlCCd0T+133mc1i4hPK/wQ6KAwrePpm5klizEYqR
ZRvbZJO5ykMjq3royeZQ69i0yOB0FMcWAJsKkxHQXOBw8sXLrFf7C3iKW9YE3JW/FuqfXVKUV2/0
l3kTqo8GUD1Bw+OtYZS6nSkT/nZnpSVcI/n6x6QhM+6q8++1eeWYqYwkdJ2CrabNKtXc2xibsZt+
IH/Pzb8yijT8yqZzvZ2VpSb2yi7ril/njL1SqGG+5J2D2u6egjDIE8auKyJKSueUZR2x3WLEkEfA
ZSm7FTi1LHbKdJ7Ug13HRyUxpAuAIgaiVlPi3fXPOsJI8KiK2lpyhVUza3KSRYM0rU000X1DF1IZ
/txTeJ1oN8H8lRYXliG9ysIQ45qOpQG3rlagFc8l5LgKrk3j+loPTX1oaPdHN+uy+I7g0PEml8uW
UTHd6hzSBDCcYJbIwdYG+cucK12tlAQc33kMhcjqFhXsOUpck1bOzIX5K4UN5EUNGbVlXa/VR+yF
Y0QAZ/FkrHvAqyxkTHq6qiGkG+NfM5M/1Lz+b5OAvA/lilCp1SXL4E1VbUWyOfFrUPNKJIJp47Ig
5bo+iADOOZB1tmy4FnhqghxvEtFvhdgCOUjCx9nPk66eU8N54FaflTRkRg1Xg9S/r38CgBQVmhbR
VciOv5FyqrqBBK2Px+4WrZ9bLZ9V8ZoQjWvCPlNWn6lQ/A5xpHZUOvP16A3D2qXMMOhD15BArugw
jAsL4quDgaE/+5b8yPV+In6eVI8lAFGZyCgRvxIQFMQjX3/UDWA5OpoXPx3lYE5NjBwIulJ5dglg
me5hE79DrIBQi47W0W3TQVbd62NXyXBAx3Iiz79Cqy8+s4OH8TDkYwb8GspDT11PXgjOlTFK8O/G
IdfUyzCDw4Tc6PtsXIIq8QqNss5rLQgDha9a831Jdjfg9zttLGiX7n2MCe/nLNG6Mqr+CaVhd3Iw
BPRxthdPhFCpKcjSLpIFUlC+3v0Pim1/W8UpQ3uG+yQM03JdmZcWkMEu5OfuqR8Tdl/YJSRwOEKa
Mv178k/5M9sQEezRYDpSODXKe4g0c3JxY9VIR+b6xQ0ByEUjIw+GA01T1QZaTTTSihncOYY1Eq42
PAtejdO5ObbvUX/lg6tpOIJ1Bv2SLBE9rDDDPRw7xSK6+r8j8OV71727OT6r/eWWnIuUq0cjWQ+/
kGPcQhsPlxxvHva9p6viNigpogdjuPIH1wrSAo6yd9oc5GZe7gr500Yw4ZH2ZJjXwiJJowMthEYg
iOZPrmBHudwYOtoqGC2yZfmbnTxBuClR8IlJU9z7vXhs/4UrhkGm4S+3ZUKFkdWHEZi6lZ6aPROp
EpP7V4Frnnkx5PHU1v1Cs565a+J/wqHQrpjOa8H2/wcBPv+edCwetMA82bhMJ7lt1kaH1b19tLoY
VnRyaDcwQg9QY6Kh1Q8nW+IYWR6ZJRSXC0F1q0RNuBqWs9HeCVRfp4ImI/mvdbGXGvPnHpdB3fgk
0qU6E3GItWe35wsJ6Ng6fiPmuT5K7ic1Qvw+E9zwddebAAPFDDDBe69AGNTR5Q30VglcmnpunioY
GrVF5lnr7aVWLobvXT+6iJn22QiCkMOHU3sSmBEXc+Gkh654uC1ZY6Fhs8FW3ko60BhCFyViLsQN
kj2qP1FVT2spaaEfD2Uf19QDm1ez4XOuU9s9nZdgv6yy3K0DP5ZVeRaTgwwLDNq/uFRTAppRh+Wq
yEzRyIMjjWjxVnBUVtmXU3DqBYzYrWh7ZR7C0/P2WOOnCue/wtdb1kOkfTlDiI+CLrVwJQFLAbbL
UM8d9KmS3zkunXpr7817vgIb8KAvjhmckigYX3fpOl3wQOBruA9R27ZHGaQVooLDf9ITXYlyW9UN
Qt87BvaoI+RVgjqjceRILZasoC+uprS3N+0kKyEELLlh+auJh1JeQN9/TEBuECOzv9d5DyExnTuO
qmQxheYUVb6U7Tefg76LLNEK/xorLyGa0ly6fgY4bpZPUPOQL4QvDabi9+pUFfMuBe07DcGJPRC2
sDepZXZ7qsk6g/CrMl87tqm3WoW0hz791K6rSnusvnVJqlXYdVLYMFdJTOTjtaX8zllWaLH7bNMj
cE2d9YH+Q+uXtVCcTPM5fC/HLQoEkLOlQVnfQ+1IcKhlzuxyVTXsMW7QbdZMby8C+mCjCrdwEuVx
NBBzSkIZWWtkNFGlU9qPHS7fFv8lZ/NN5pWqCuuwHJD2afmj000uZ/lBxO9lsSBwQ5a+WuFyA06D
2affwAjpG6q0mT3DEna19wSuikjU1xQ5EBv2i1NRUso5CgUogaYUxlRdFQfAqIySof9pZL/Tp/2M
W8iWbi5YI69vMK69kbfNlVVzpjySqeglSgsD/9E0Lz+0wae8QaJVehX+CqN9Hibmcc7ELP/A/8ob
ragbWL7vTNxHdo8SMtzZTzCTnqD3GzIZe2LHy3M4dBDEi3mqBm+nOHvdEu2F1WM06tzuBEyR2Ndt
ip9S9/Da2piCSuUkVDhwiI0udv+qnFwQfRWxulQs1hKxpOeHjQzFE+ZGCi1KseduC/uNNfpmz+At
rvjfsOXUmuss6QWHqvKW9OTjorLQQsS0Q+ph3pfn3Ck5gj2fIg8dcqeiCC0YZ7Gd/cMqwjLh5Nc6
BtI4j32cXNYoWCEiYVOjR9nWx/u5W4iGropMQocSSti63K7BZsN5BHPo2EYVWwq92yjzuL3XZwCu
j6PW3uLZubDr1omUblSWEO4JjWoBvx6QMtS+4KJ8iZAMg0SAskwAoey2KuM1VazP68QJur+edJt3
nAqXr8gJYpfh3D4Z/lJ6MiGww0MDLr9B35r8mhef2256mFhQrcdqAktbKgPcWbnD03vxjnnYO+QI
R1vtluGD2A8lfpFqxFCwUGvgR3WHZXZ31A/cuX7z9BRPidTU326aZ807DKMJNTdmW4S56pszu7aD
ruaLxIMP7X6Mf0GC9N4WzjU4SEGkofnfRGN3Xzrlkq9C7MBsyL3nd3aZFSRtz+u5vkzykoAFiLWj
BpNS5KgFdl8aqjqZ45igSQc1hzhakB5SQgLgthAAW2xWDxN5MLX10SIk6sCSOr9MMM7NY1Bb46fy
oDoHbNrGjzkB60t8aeOtcHCt0tAr8D8i/o8kRsxkQscxNbPa8azkPlcrwz9gMvG/Zcvvxj+Zq07K
jLS6iWLQjVpURdS1QBmyetsAeUQUSF/Yk1lWSdzl7Y2p7bpOD6ZAowhOn91WVGcFblL7vojxZ9I8
0F66W812fbBQuxeFVGaO/VF9OzP2wSRjlNB1svqAyOFPCWHuZz7wY1Ktm1GMJNuJ7jx2ovzIPqoZ
WwXrr/hUcJpBwkcOdxl6LlyfTjopiGQTAYvlP6YBkKE2DegB6bGRyyy+z4kdk/tL9vCQJ6Dhcmwa
6xayBrqhE+QdRrdPNbTWM/NfTdkMkzOcxG27gcPElD7GA7zE5y73Fstc5havtZMu0S8aUWYJWwwd
TL9fOd08+gD7DOPmI+FiiGT6DTnoG9j6gGyTRArY5ZAzxLBUrhjd7+Ldj+aKJidlkfPiEwSb/BfC
DBEYMyFyqcjU5P3ZmDYuSjTGesVtWhHsm4cpmWkBrnFkJ1aXrWyemjJu+/jI1CHOUP5AxX0pvi/1
WmRgw1AbUK5ZrFdOuekNWsatPMq4lp2R12/B9FAMQji1KkGJDTJX8/Y1+fIuoPSrCpb8uDoJfIcI
rYvP6p8SojTtyCKO6J3oDLtzMXOG7tIYxYUkyFWVr2RgmcvP0sUplcZCISa32ng/TanoAuacWe7M
2ZhBel7Z/xlMbXJ+4R1RUAZL9HBgUfU6ziVqBzPKRhTWda1NtRsJbD8/IVrw2PCsXWRGq9WZZ5Ja
WoVsCAwBJmyGW/+DLrtTmNPnV4YSs/Rv6txthTzoB1d9dlgUHybOtL9I6mvN9gKUFxaaCLfZScJr
mWWLDDsEiPALvXfzJKXmaUjhl5AaHyos8gDLv9xRxnHzXaH9yv7uwIvnOVXRVY5/0pHE/MQSenkk
tEKqNMxGJVgDXw26bNoEx9cwek54Jc/lARiI7F4Vo8P7kmXz8qu8h3YaiWwDhYTACMAZKLHHu+JB
wMD7ROQyIDmCj79YoEbR6nSWWCk8uKwC4dDTSPZL6smvbe4qd5AW7+WrDp5PY1lEaJXjep92XT4o
u/kDjCYw8ILde2noZDgPKA1onknD7aNq1tYgje1Elsw6AXXbnk1ZkwUeO4FXEslVsOJB8w28SEQI
C+S6pfmym5oz/k4V1gwrOBaQlwb0f9RyRA/9XsYSsGl09HC7rcfYyk7Aazbfh6E6rCSd2WMOIVRD
xz3WyTn6JJW1D1v/UQ8Lx1Y+hG/F9BGHAHjc4hf1/yjQjBctZU5LWyHx1s5BRO4rckpPtxtU+1sf
l1aPnMrIPVk3pMHm/xKKVqbeHF1v2Pqio3r0cAMMQOUI58mxCO1tN6AShhJxzUYan52WKxQcBZWw
VZmxkCutq77TeRpHqVa+M3IOcpDqK7k7nJnejSYq0lrRM9e5dZaYT1DfacAouep6/LPxmc62tqLy
S7QvZOitFVD8G6lxozziDNWe4Lmpn6zRr/8GOsa8n9mnfr7z7hBl7P+u3+xnTrs0H9XcfgQr3NYH
bq0qccU5aCwouIfaA1VyT9akYdRHbV6z/poZpc9+6Z2OrmER1EKa3hSr/nD2aHT3XTwNmC4cZ/7E
rtqIBgyyo/SG92d3d1/a4sXq7ZBGcNcLm0h5gaOrSUiA25LPHBz6N5M5jaBW3VLkYvw4ttffaX+b
d/26fvZ0i9Vjhy/k7nHz9ezLIkSjIQrnc1KmFn4jWNRwe0f3GqAc6Px3elKzIqnRhs5dM2bhDGZK
psXgurunvz6KGnsL8F2wIDPMOtNx4oafjMXjgZiOF8lwgeqjtRY2C+S5wFLdrRZG/b0IYZklYCBi
4xfS8OBVJXpd/MxtSM2WUMP0atmP4oeqZiS0NKAF+U1SapUXWBh1WlLLcWyeqtmrwVdzuurd1zqa
dd2YcuAGvwwV+7Ubjmw0WwXQiuI9BQl/Fdo4liuDb8e8y2Rxkspy07JVymj1v4hi9om7WnW422fh
LamrDDceMbamlfmDK/aqDE9brl2EyU9/Y/CjHFZ6aShPUQkv488qjEPO1wARKt1zjNsLDpNbpTro
r8f/gfpsbOoFsVCxzMTTbXUBLlhufUzgnPpC1r/DCyghsn+clp5d3nIfkJYTItkZUAUOHUVcMsPT
EIblX8iPaWJd5ikQ5IsfPY4+1XvX8fSHGpd/qseMN6YmAUEoWUpx5TnqJXokv2mDZHZ9ikmtVMmH
MVIacfDJHma2HrDpdMGo3gm9AqrcaEsGG2yIHKrt6gjYKfOrvumIsWUg7CB/akF7nQVHTYzVspvu
TgpXX/ZWnqmVq9Yfg14eKiFAbsWqrDDkMc+J6yYX5NhdmuLQyvIQVVqTrZjDXjETrMWbqucVuApd
paB5QUrMXnmhim5ujQr+1eIGYS53zPxlaHH4pglW3tEIoWy5UV032az/l7lD9nF80RiRvvc3pF43
uOTJZlcUWoZylH8uiOTILV4AvzH9JvaHlz5udZ1xrX9E0hJ2/xCOpgUFos6+dUJK+CRe++U4qzsb
fidTLd2eLpQNUSMA4IC4v4LxLD8FVXCvknIOdUdsnWCax+Dqr0tmZtC5DVCrd6g1pr1faAWoWh55
YQ/sovTeHv+4Ey1J5N0k30gCEoJKqVeZVIn3aeF/FTR/wpx3TR5eKaG6AGmzyOfEM+Qg8g4V3jM1
Ju+ERwPKwg0R/hE7LwKtjmZNPZuBzIx/sAr//8kj1r9EbtDThPexdk3/Xga8nAX5iLr+KBIDaBa5
xWe0EDlQ0jpxWFbgeu6T9B5rjmLX3m3REoy7tai8vKXg5VBbIRzCZ4+bDqxC420XcSx6Uex58ZYP
gOhzFbWSbk9XtYzBhycWO9HntMPl8xvIU06UMeXrDGwesm8mJXxULKbBS9sEIZvygpinsFJyamVl
4+utyPUmkHfVeV5MwalApnZHpo4fZgBwhG6vJ6TRVC2hGTYfpaQlvXaNwIM19XbH3956PcFidxyW
2l0gMkj1foQtK00iOy8EPGv5rOTmApQHxKld/+E4TSJ8WVMtZNBzWyyv0KalaDpndbsYqA3nT06T
JkOuRbgwDc1mNk/LPTE7gJjZaorGPOB3rgb4/WDyL1JLIxDAyQqqkD+/eTR/cisLRRbTBAhKCQ68
2N5K/Scm7jFudIN0DXLAJJmMOiw+ZeT1w2YV6ZPfriqbJZg2xyUuNHLT4hKD96NNbatgb5Ur8zMR
1twutiTo9gCDe9aRtM3tU0eQHs9NouwOxQoI2PaiFYBS1kt86AHJfJTnFlpRAwsjM1glGSffc8Xd
ciBipcxxfAsZ7EkFY4Y7LP5ZsBZo5gh7aedm6P+lC1L6IcbrFHk2OgONUgtXvza+iR46pTmpsVfR
Iri2ZnNOFDNBRx9SuHqku0/KBkpTStf9ZV/+DKo6ynZtmD5HlUW67H/NpKltROJYSTxNhAAG3lLL
fEHXxHz2EqEuhk2daTCbHXbYf5p83ufJa+kszor2bMETOEaGF4jzT1NAOov7jm87he/7yqJIojCc
UsmxmOciAnfsuWYRG22/l081itH1LVl96fx2rcyKBdIdpPdmiyxQfRdM9yxGTF9BQsE5H9kRJCos
HvD0K8WEwicf1RilhvWAWfqZj9ZvKZxOLUqPbdgORIQkViuAgS+x1+v1C7JPRfWirG08cStURZMl
JqsbvesBQE6T+AoQfxWlKPFZJofe+ROmpmbCtK4CnhAyqqoznjw94Tjs/jiZfBY8fORu+hxuu3Kf
VKoU7qnyLxt679kEaMIFy4yLie1awdh5u0Xe8jQT+DUgfzxT+4Vs9opACU/iKxDnSjaHn/pBB74D
fvlQPanPyhY3uUYgq5an1beX8cUegCxrYTCsU8n9M4Vi0dRgG0BavQOF73ZJ+ie7egg53UNWICfi
MSYPx0sFxG/XIzMDhvdT4oD54rovcau6CmMQ+EMZzz84V3R7rf+CKj9r5Iozu7BvZuL83UfTyPaA
6D0H3og/ZYEQhW72P3TcTKY8K505Zzdh39pWx7qCwY1rT0hy6QkV02BaSoLvRybd3llROOlLzgjG
0+BlHNLtl7eITpaWZGfEUTm4d4J7/+IJ2pjLrKOck8pQmO49Y54f9ziB09TgQyMVk50H7mF+kEUP
Vcz9R0QkcbwAC9P4OJQ7xYwXXyYSWMaIsTq/6GcZCKR7WfppgsAIbzUBCHmy7YyVHhmMwmqCkLm9
OPmjbH/FOXdyvWuwNdFKJIMTW8XaAGNHNcGWJPKwvFnZZ/dx2qzPkF2EEj0ulFqQ4v0OM/GcCqZa
ogaprSkTzIEVBHL2R49IFoSHUInORF7n1V+1I+GEsBj2d5jU2zfPBc99WHhPZqoa6zU9nW51vpUm
ReOIsWB5Rg5PA1tPN0owFlJg9zMGm0vTOChyIVSWJxQlLEfHqrzJmfddlalrt9BmEgHPpWH2BqA2
r34N9t/fgOf9tD1rBYgib6WrVAWFYo8JgFkWfgtQnWdn68yAD8bYx1PcfpIaut0X3Y9B6I6jr836
xzErIrVj11TqpuFqqqcEe2IUjnxxG9wlU08yTRB1EyoBuqU/v/eCYVOJBwwVjt/1vQSRfe9XGiac
snP2+1zMESBUqHtwQXmWHWOyPwoT9pvEgTU6cfQJoKWpAgIIR2mgTyJsvrarNS0owVysqSZtK353
Cq9KwH/ZpsFzmLaLoYDKFaZFnlFAA98z9axALt5zXKGV1dT9eH5eWKpSGujPSzdkI46K40TbT8tE
bZqYuGHGM8Iw4jjFdW9hPKgLNh1Y+0yRwHxXK7xmCaI8cckJ1klgzhBihRKkxRi+wGbG3/GbkBfK
XWF+YrGK2yHF4kl5bqYBobHywUd3kb6ZJ6Vc2DFn7eOrgoR+8bxI8Esz8J1DYpjNDX2+WrwyJ6gP
nE6jyCPPZphzGa8GWst95tV4hgpF5MXHDEoxbETLSOFJAIh0RNxYOfn8oW6HjhJOlc0avHDlrqpI
eDINPN9AKBxqaitzUhPDwya/j61+2qUilENOC8jrSOuQzJonTQcIdR4AIqUzSH1RqOkhjyOm9B0x
BMcFFFQAEl00/3Ib1avIQWhiCUjPj+eJniW0bYxIYAj1lJN9UWnS9sImEGmtLGgvSRT08w7sCY81
qgEPDnxT3wAnj6YNVwbA06CFadk9QJntqvlOHWVnucyLgsFekbpv6c/kYCJNRWCBhgicTcHXbj5/
4E5VWCVVYREvuQ5Vd726amkBp66IPvsoa7XCSbKD+tVU6S/GC6CupMb6DWE8aMwetBZEBxuEU4YF
24FcvvjqDI+aOm3Bf8tw0c+N6Yyx70Uhw147Qip+JraRAWuEbWjAPlNvqEK46/DPoOx/viCiiqSs
bCBt7eoT1GB4PCDo69vP0Gfb2TxeZsdzdBc4bjNiA5B9qTBnGxSOSviERU0cROUKm4c4i2MpYLNY
LficUai/iBzLkNWt2TcXHTP0z/ykYe99OCM7632yZMKWlrl2xRW6vu0fkhggG82Bwln/6tTDZQPb
Iph46p2VPl6Z6A+or9Wgpuz1wj8KMc45fyi2q6S5fZ++gep8z5FHFV4mYzsnR55kJF4YW4rrZe6N
cVBtqmqfD1qLjBpM6253z0IV8CwISQlAJh8UZCEClCc4a7ayrj3h1r7k/GzHQDqO59dK/F9cfVz0
pq1QMLa4YgVAQkaXxKmy1L7c+IRcwAxmbZXZV277KxK0BCUI6KaZkWiAGN2sb4y5BjnpiJ7qLfjF
N5N3EqTn05ejjUmWftXGyZsrT+QLJ7rBz/NWQqsXWr+XspSKMvQHDnMSN6fOMLHtUfF737dQn5Ob
Pavr1Nqb1ErXGCOvsGjbCAuwpySWHb4iD2J5abWV4peejwjNziPBYDvD5HX9GKuPd90CRG1O1xkv
Xfa6iL0AH1rKJX7mYCRBlEKBYQ1FN6W6v6dkjgvO6C4PlOVmNQIXMd53+gDeJ4+awGHPhvT4sxp/
kXp0LHR4oaMr4nSmZYDLeFhqY7BmhywxfEdYlEi4wtC1f2vqcAq7jvpEvCL+86sDYKwJrXPIxu62
GxmpwvFJfq/RtZiFXqwZRVmR/izQZuvU5DDZjLC8TD7GPxOnoT8DpedgqK25QVNXCAe1gtDRXNiR
WCTVgPRLi7d+tcXLSw3XnecXCE49gLNMb/48aAmTGl8HzwUjJLsF2f/jIK4dlMD4O/R3KVaDNvUs
4uYVbi1pXT4VRRtty3/5QWSZwz7J1+c2gluanK9pq67u4fMX7dR+fvJIjRF+MOrwGK++KbxfLSvl
jcxyx5mcIXo3hoL3fpy3yq5ce/2HUOXrFRICA7iWKv/NelgSvFrXJFrjeQ5nLBpa7+jbSfBzrUgl
FU2J3Rse7I/sQaYy4ZbQbuLGlUC5HRvJ24uePLSwKh80ucSlEQLNLa+Px7ujh8hQ4mjNEghxjNwJ
fVpGe3PkPzGMj5+YbbtE10IDsXu+U0YoRWVtJuzsh89F4tDGEg2niFcbgrVZqNcPwmC8EwchrYpv
OCHuP64ebK3q3ej6oF9rAHpfDUgOAULIVRifeVTGPB+eBFOtoCB/qE9eMVjzU+xKCEJJqNtkhlzN
QWuVIhjyNR6E41vNNCf6Hwin8eOt3VG+wO/vaBVoc6T9lX+hPQTkHksHq4SPPKzn7DMe3PXbJD2h
0QuMKsTY1iUUM06FK6+9E6xpfIZqTEfplCPXl6bYB4/sCARIPW2pazpDLGoEwcJ10u1Ic1VSWBZ0
eo0wZ4XMF5wJof54H/9K32LsI3AQLw2D7BmxfvEUS3oNIMWCT8flWh0bsd2ABbzbdWY6840sA3Fe
WJ1HJdfb0NC8auSsxEz2B/7gcGOfxaCIR3UDjK9p7Q0PpmOcaYaKaQ0IRbUaOCxrfIDBOaubwNQd
MRIJV7jeJcDGvoWmgXmwVQf7QagIrPQEkSFIZZhow+SMyBpIEFJ2M2a42h4T1UBW2mfBxAQJppU+
HWHZKbMDP7zXWZAJQIrcqCFkf1y0M4zA00Fe5DRHpG4u+Li/FHfxedXQAi/+8lrB1basF6+HSBFp
J4AFx37F8ED4oitt318VQQUlvmBGuX+81tCo7JFcDClohWfBujcH1Gt7SgGjpIDpelddF5JtliPW
h1nL8nwImTzx0wnaB5C8pOYpiWbyo9LJwG57XB8LZ5XZJXyNDdjRs3IccuG+H/PbmqFEJh+zi0fx
4V8b3XhbmlEIizLM/TjQJNisWQv7LZ8bMaq9pvmF+hSAG74evFPaUIVn6SIHfze0cnZ06oe7iT9j
5jCIDSsj9vjE1CI6MPpvCh5BFPjPs4bzrJtfRtXlx6KGHEAzXQqOogy2gP5Ni0xwmEmkkB0OXFRJ
p4ueLxdiJXyE6yaKCHxDhElBFGOASbhOceSVS8DXBNKmeYtWjvGMWWhmNIovjZv7MhYb2kYGhWX3
biRh4h5enC0K1HghjyPyqgAzJv4S/K78NbiPaS9JYhStij7uRWwvXRkXhjn0BOQ1e6Oisg5yiv1L
pjHKeZ7ljxkSmrfHpgywVAdEjCWUv4jRRMSwRQ02gMoP0cVVvdqOZQVPqsKiYXikKwHrIoHsXzUv
D3sNcV3kTxCC1R54yS7K+qCF7wVkdw82jiSsZaP13QJXTNQqWtCDROsh59XhAL6OlvgGaGWYB5bJ
H9DCQh2mMrzpk01chUeNmOKzy8gvYmsv963m+/CJbhgb/ZO5M257+3EIq+vFFDTUQO9pgrACT9vM
jamwKFOgGsdZvhFNbPG8NxYhoU78iI4U3w4G65daTY/Q7OvViZqyVgn150iiWitZBjZWHChmuRDK
gtuSO96e/QY1tHxbnhSQUf4aHjxXBHoR9lhKg8PjxUGXTqefzmuHcEvxwiqNV9Gsc0cd1iB+xaBC
YdgYm0ogQVVcT8hFKQBkEJzBBmlEiSZmvvBo60/RmJd3ej8CIsZdc92KymQUlgfBuf+66X3F7AL9
6cZKqTr6YHywx2PrKi6XxHbjvM2XOMD5USI3kQd+w2ZArDOcH4iSbyotTNOBYTVUiuzNhhEg5Lbx
e1+QDXWiP2uOYPxnWchmep3Ncu8ChGdjYAspoaow6aKnrNWQ6cbY+LzHk2enzi5uw7RZ62UtwirZ
7nbD0srd015WuBZ9NiHX5E3uM2xjkob+ltJrygbxNZTUJXxqkPtWrStnITKtrYSV2vUkdVz9/T3r
K4MQDTySGIPiDquAdRyXpGiRwdTs/IvEwr6drvwr8xBTfrusOtaSpi/8jyy+JfA1MgjJ5P2a2WT2
klsSFUkD9+VoM4HBg94aKW5yb0n7XXkabJTqXNe3Wi8Q8l6pn3OzSkcosC6F2CVD+jUCamC3a7sN
VGz2+vLEoO2pTIXxKGidN+XniiIFY+AlpJkOpZUFCeG6A6MK+VGWFfnCvtIGA8f2+VaU6bBTf9tG
qDrS19yvlagx9ZMlDt/CFG9U1telNlD+Q1VWdO0vR1enDvzMFfpyAtbyQG8d/e30KIYGvBmpG1fT
xAmVbyu2uX4X/ZogG9M8rxirvehk7kS5gPMQmZMPk+4+5UdDajpb3o/C/6ciUXwjRSZM8damCbZW
7t+EbGL1nHi9lx1pCxRFXesixGkFz4GvXf3uHz6gEucgVKhqRhw2/6co/eLDPQwyScE0yEfstjyQ
rbwE7/nY7PO6Owo9G8SZ03uMiXSvUEtwB6958hm+5HxOh2cSL2H2Bs9ADE7SGkvhlTjjlUQVqo4y
DMjwADrm82ZeFvQMysByG1xO+y6CQboEscC2gxci85p7Xmpqkjx+zXDlFJM9p5AtphGnB4BkpO9s
VguohtUFBw8gQ6lDOoomdkFsXs6/LXJYcHAhixxB8kzh+dph7/CtrqjtenTVseDgzjUzcXyhTKO/
Dm1YGlbDvxvkRvwnDef7Uq/VAQEONovwqc791nelycmh87HQzKGT7HOwNGJWRe0tYlHZ4OjFrRQZ
sMbNKaGV6N1qUgwmbLaiPN8C3q9eYoUekF7O4dO1FvJal55Uuqch+4nk69ILzqKQAP73M6rrwg25
HnVEjue3O24oQDFVOO/1NuUUVsvf+NzTt92XBua5aqDD1GORB+l56btdRvAyw4emgoVjRDykr0WX
lw2I6Wt8d9T4/a+Jl3+N2bwv8aAfBbuKX+fgwIIfnLP1HlCRxT6yZgWhrZY8l8wL2DIdbQRGf4Zb
Uu9B80ULpQ6ZDDrHDr7ebR1VNqHJfik63J693IG+VK5tahD504WkCsuOWYy1H5WqxaWYV1t6Cln5
aGR9L6pdHGDcyqU78tmPvSfJ+EIat02dYNA+ccChFge5eQHE6guBCxOPw5UHeZGLUj7HU5Q1UH2o
KWKp1/2LptC6XYb0L/cGHXLupVMjcbrJinJ1HAOV2ayMl9Xjgp8piiiWQOydhFHPqTaEPOjpGdZI
Q+A7IsqmK+tPm+iqOdtXRuT8KqrEj9f1ASUlL4YiNj0Mkv/UqUDUN9LIzGiu6e6u7wPXHZNvAL+r
UqE5Yot1t2JiSRMlJmbbJJjsdY4v67n8d6Ua7X+xJIbuKgTkzZ3yOLMdFxQfMLoHlWu9I7v3D1lE
Cd52kqcYW9xNcQznKZUPyphrzIlPOQvg+nNcXN7x2vz1Wz0dgr+CTlEpawSnr28nasPFwM+ltXMl
Mu37/PrWWFGuskYGYFvwG8RX5L1jEhS1nx5ZxUoz756RkbARUWuNwlFVdOTozD7pavcmLzU4/gXa
GqR8OYvdQySQT0dqE2yVVoycS4AmLKbTCHY/bACe1eJYwDntENNlxgkUEOf/CqFNBm5f3/JGC3b6
OySNDlJKPzpp1g2Ol7MEjBILkaLLhVU8La+LrQqLHdMY0mZ41ta5F//4MhV2upWAZhdQlSXsXHrb
pX4P0bysaeQWoYkfBgy6Dc8tzFhQ+X3dNvzulf4c4We7glTS8nqTEKv90saCZ5EXsRZxDEBoHWk6
5huk9tEagTue5+4UnF7t4SNScs9kCeB04QO0UBwVOtODXuBKy2/BcCWOCn3IeeT01iHxyZci5+3m
Q7I4HzrLTx4Bz/4QrxNnbUuqA51baRptXUeF7yDkDcuknhExUMJhBsY2cEQfxkB0zek82hVfSnsk
ZEqtkGR7Fcc0JrOgWJ677gzDPXuOA3iam8Kj1Lbu2tLYItthCEBFNZrGdbSbmDBgrJGEcAkkH30W
i8N3h5AuhXxRpxwe/OuYmXCoBMxk0n71Z9DdhqaXCsityrjmKixYj0FH/A0GYXQZTanIr5J5x6Bt
XCThZEM7B7xiZ/YCYbNQpXa0aos5gkVwQK42asGjuugYbWkzBUQOysICFCD9UN8ulsgSmku5ieh9
1emaY9kXvqPeYGOqpR23kmcAIl4SCzAQ9zmPaXLgfVfma5sjH+c/6+5NLVj70sjKzEiJ9hIBk7EX
U7x3QAeNWtboPEyMKwxmNm1L4Vtz606O3v6gcLgdZ825Ln+bhrcItG/laL4wm7x2mUvlaXUdfikI
avJk/y2dIVCxvHKFdbOf2mFm87ahpinUJRFMyCP6o0tx5FLwY71jyIyweSpQk099TBDTNn9pDfdq
W+sAwodYNHWSdIyEPx1Pyf7H+fjWYxbTvNqBpEuvw321zPxYBsgT2239E3PpqsQ/ve7uGxMdYBIg
h5j48kfhB8oML4whk6abNDV1cgiGFBtwqWxozjjlsjnEtjya9ILf9yMiL9jjGmZbjYIAOWibANH8
vcFhFdQjcIB44lb2QcxDbOx0711AdwZDI5TU43D2byhMNIe2M6RXub2ZTSQUswiN/vdPx7DedzFB
+N52rM5ZVadxMnC12Ewr/jX9yaEcaT1HbCe8/1o0q6bUNE7ZWKN+jTZi4n5WFU3F8T5M5TBy23l3
UAbhmH/9ka933RTzSfIAzEoocQzh1+8al7jwMZSBqD1TDYkzslQ2h4d9F/Gb+TwqayBOxH00dpRS
Ya7aYYD6sk8xEoIsxbkjbFPYnQUV4VdRlmPQyGneo2FDtCJCbboU+nN2O+vEIVKRpH0FnuA1OchM
s8ZuMdFZWTYnmzhEaebRA8AGI9d2jS5a0h7Oq6anW2cL/pm+Z3Cvcz1V0TQwcB294xm0p0EL2g53
NBxdCQY+bpu9DaPgICCYVtO469IjIQddpoQ0cgNCfT+JVVM46vHp4hmO9DwVIazLmhxSN3IhAXhI
SCA7bVh+KDN+SOLz86K6SNswXcr7DbOGST8LFceLwlzN9sLmill/lctnl919fV+eEENe42VuxErY
/xmOIOVw3/dMIUeFi69pBNcpA8ILqRPlPSu7CwSDqFG3bXc2TW50URw9tmBudHJ1YBgoFYuq3h8U
E2vLohNnkLv4EziW5wiNyZLUnKPn70t14RoszYChjn/0Ej27oDDtzTRTo1wDKi7CbCYs0/QX3sLk
/duze8m+Gxrm6wcugZIh2JjYzpAkJbc6nvB1ktt7b1Pmo7bhBGAoHkBxAsGHdB2HXzpSON9V6x4C
T0H2SKB7T8KvJ3FU5GMRwXIOBDJLnthwtWlnA2eRCztp+1iSHOGPJ4Rc+BMMqDBrRMPedVMaFjWL
fr/zj7jFc3fKTNEY94BHezEC9uG9IeNuIy/IseUESHeynkskt9Snf+MFIv0wDck1FWz9umdxXiif
vBM1Mq/7YfTE5dVoHidQLhlGJlk7uFD85RsLogYL2LBps2uq3Fldh8UYFIY49LNEqEBWSSWZLcKQ
ZB7pWPz4sC2P7spr826l8shVIdqMTxMm2FduXZ7V5sYit/NeCqDh7A6kB4/i7Q+ei29wGGi0o45D
PZRkQ3lRdIsbTmJGj4CSqOjbcd0+4WPYYQTGVGcddlrPEymU+z9vj8iNCNo+KNbtBJhETQ0LFCZC
X58dL6KHKRspqxGOVBagKV1P4piWtvjjWZC6x85utFa/sZkv/1tBkXtWl8hxL1pLwMQZCFhyhIkH
3oDot5qkZ7VeuAjZrN6bK56QG9CwkTvHef/ju/uf2k21GbFBcCt7UgUmLfjLKeIhKL6OgoA5kOa/
1vjElwq1icjjQkDJNQ2Cf6P4A0083XAgPe2+YCk3QFKg42f1BmfxJoJoCKXI0LVd7Jca1DzW8wDU
5MVhmALFju/64xcXlqBrXM4aBVv/P5gbEI6T13NIvKMbe62Chl6BbcfARY2yCiyL1ulCZ26YixIp
bNUp1Ac+QoF+hhtaWcnRRzvkCEH/eucao82AXJIiMrIonZ+9a5/Yi9hJPxbzR3t6N9koFzOpy+58
pPbr9/rEtCTt7F/kGoy9VyxjWe6W3Gsr93sCl8kqhTr5D2V5OotMR+GdlYPdCUB49S6gTcSlGP8y
JW0gGW01RNBG/LFv6QN4qg3n6llI943pa5mlk0ptJ3P+IGVLA4wQp23T5yMl4cSgLfy2lTA+O5JT
s212nBXgS6yuSJP4N+yLlm6lnXKIz5ehDx2RsTfd/RRChNFCQ9vAklr4BgPBb8oJbuVWKBZ8WwvK
TP8yMyHWJPINOLPIZOJMSndo0SK4BrjVFt0HdTLyyS6Ng+p5MrWGXK+zx25682wG1s6NJqsBcSSW
0uFJYSW5f6Ksrovun37WUUFlU6JWvpDHhRwUF8APKqDmWXA/SNSW6GDO9QLcnqyLRzh4Y0BKM2Hp
OwRiBS82Mha8o3nB5f2AgG3IUVFWcTq//Ta86daXvjr9ScurBFB4TuhRvY8G9tpXk/oPBtLecokS
/tAw2arun3OwamY435UyHqErMhZqq1flsByMncWBfvnhA/Hqjwv6oit1T2O4TgobWhuszynO9wpj
ZNl1JfgdjrBnX8ylJd1IvxQ0oUA8Y0I/xmSpVoV+LsAQr6tGdXNtW/f9hO2qaU2asOEmOyhhY/LP
dJ2TrS+XIOrt3fpQ8Ex7zwynUFzYxAqzAd0GkVtsbUES6FZgBb4t6ZcPnBTInEhrASFfYwnPas+h
TVyoRDy1a2zSqxoeGc9bakPaWWFAfybNAE8cYSr4pcyLG/dSOuAPQSSHRejc3YijA5z8BnnjRdR6
AKwfLfEkvdqrDBLDYACcBN35BRSdfo0H6zfC9msZ4EtxlR1jewgbcqQxN92bWSbe7gby4jLXSj1W
Gf5RumpUzEpGEBYdJFPiW4AlZ/seCbHB8g1Wmrt9ilzewGD3rZd7UC1waXwQJwHbKKqJQqIYEIRL
LrUUqLzlWWrOsRvLQgRTU8+b2v/MZs2In2JZYgPMortXLWfuMV2BOfREv+iF9CN7LvVfyEzxdBH7
sZEViOC/is9QUx5NvTUiShslcvWrs7GvsbnLatuQFnp4mOgGZ2zBdog90GvzmCLOaFSa+vZBty5+
i9+5Cy7De4ko9mxGwL3kslz1Dp5Ghcv3wFi9IbclHWwC7AZlIDn+xVevtv8q6K4rC3bwugiZQl84
/vOSXaJAQqh2mBAmCv7V5IzhFN2w1Y1bwpMVy1ur04GP123Dbdf999NH0Ff09NWYcD4bsyxYrWFi
J2T5HnL+76xLfvp91QGDk8rLudLXQP7SJ2OuPDSw85vvZoQgB/y6c9+WbPbo0wcWmeWGYXY5z+6j
oiNLiKf+GFRL6nzRi+UE6NBGkKvFLVdVB++RUMzQSTpi+oM17xGpaVI6oAxqAQ5Rsk5CuFTpuCmX
pbRpEvzVXH+BqXFfwsKZyE33SapqxsFCicywEm7hdyqpZqJ1DxhEvOCdbrjWuh8H4BGbnQlce7f3
QWa8mIX/cVxUdLoZmoHp6O8hnBNbz+46ufeqXJvpEUFvNdT7IAAdbkhwy3cyhe78vUjL3pWb23uT
uUWkGF+ZMS2GbcfPkpGtyPPbLZUaodP1x1E2Iu1yRmvz6PB6zl7ryOK/K0t66XNDKsApgfvy5GUg
kV+ZxACqUcweUkb2RCLbzA58hQd5Bk0s4rWUV+JvA5/3R0anBpVrLD4316Y3z/vYn0t9iyNJarHX
wQHiA9XEUZskD10Vg7U4B3qGAjYoNjVJRpnYx13ua6zd5ueZ7DbEML1r0iP3Hr7T9oGum+OWYynN
rnUkoiz0fOdJjY9aadUCIFFwFJO3Ts+Ju02kxMhfMqh+Fl0WZg26e6k+ox/ZbfVtZXlVFuj5DAys
setr7qhSgDujdN8QrTr9bwJTHeivRDZPC4XzLrDlOYakPtzuMbb+Msomd2Eor0AlmE59g28395yN
zGbIf58l+3oQjzjdFkBco+4TwU0dhuM1htibqSPX2sYwmYvCevvw7Fs4OjQ/mYMfYb42niGbBOT2
ztej0RusduJDZBloYSytpvpXHCM8DsKgOPfywNrxkMy5JlYM7LgTRTwxkmh2jr64OakwIQ8sh7x8
lIwqV6pYFk4+RsRCrC9mT992w0wOaAAkFI/WksiIcIaPxeMiQqv/+aKQz+N07jwGi2zlsw7xuZYc
wcWdocatDPwqjp4Rh+4LTfpBxbQY64yznp+WP+QLYsXWrnNVyek64Q2O8WvmRiVrgKxfdvXIMWMz
Nw2P1CF+CtLbXD8bmmNIfWSvt3ULcmNA4Qd3TQU2iPOte/3yt2eEWlASiKFY/5TUn2SaXEG+fUki
1O9PmuRSjl96pVvtUxyeyNFp45VnLYx7aab6AcnkT11ns1QCL2Tu78DPVeP0Xi+iDxRLUoigU67v
DMQvyHtD2r6LiyqqJ4TKSHB8HclKwLNUua4kiuvuLzGdynu6CzHqzG6ShJeZ9MYyMQrcckYNaVXN
axrX9q+AmexgFK8+jAKFy+wOxLWEDolzIk3l+raT3pZo5xcGtlHnxUw8K6cxly+JWms3EBh2cNyB
ATOKB/aoFAbiJIalTjDyZLPQwOB3MOiPb2AQ+X6v5XNSYY/qLdG4VsvOwJHizjtA7Jt3E0Hhpykk
ErUonjpjSApm8s0x8AHB94wJ1STjP/C5WdGvBURPqAyJCm/zoU9RWFdwtgnszFJhcttenSu77GnZ
8OYl4m/zQ/w0Mx8aPP3yPHWNUQgyemNYJZg98xfxjYSOJ4LCZf1v4BW+hspRmRtYbnlxT9nX7HmY
nSnZWatkW0lAkgXA11KCzT2ViSbm+jQ/L10Bht9r4o3Fb/byfu+t/JvjyCftyvj2C/wvPWJt1h3i
9pwNldezXDZ4R8nXrwKLdi7Hfy/Vr98gv9SkgJwO3QSBueDHIIpI/XlbGJhkSGQN2Fh+2QmYZ1/1
3BX0FhVqxNgKEe41wM6zBBAAUMbJItJehvwclBfQJJOGzqQb5e1ftFZQbjiHtxvmd0vugzHiF1IM
+YnNrZpyPfCnimDMzfWvN1guBUzSIKrgT/0GP3OJgAoH9h79GtHciE8BqWmQ6vRXVc58UW9D/KJO
Lru8BlaaQ0G4LFEvLD+UDVy6Fji2nwsnxl4dSvdcai+lc/4vyxt1WDOeKvQmTj/Mk8pWyhq77FK2
go1To0pBntzSnY63LlLEDzfNq7o6PnazB0HrOCPhqYjXq19N3R3rNMmgybTBARsGxzStUl6SaC0j
nxe6mWgTQxCT/2L98sDEeQeBZ1yWOyMpse6ehBRwfahtJn2JVpm3I6XjglECVECpo0lBZkTEmXLs
AIiR+kVIJFoMpvwhbpBqq6uVxmOnZSqY0efzeGnVqyC9xITvILZmvStH4NYDrbgT+knRV2d5FpS8
+SaZ+fxV4Wk8XrCW1xW3PYZF9DYIWXuS8P/Cy/HqaTwtd9Mqb2QUzr5zG0NUxUkYfAUTQ0ogY5Eu
lQ0reqs2i9h/QCLcsEYqhgq8m7A/tncO5asaTgeZOQluttjILOYUXEP4bFzdo5raoXkbY1ev4mSO
Kk+SK0Gnz9s55iyWllol1aEf1hAXzOTN2U1++Kf4jkngD8H9K2HrYg3BX7FoxZ0HhgWeW3kczPeq
jRpYzYdXzZd62k0yfrIO0t1WPthkUF1oEF55Ov5MS7OMtO6CwlyiWdFamWIrqWtGko5izKpmOIb9
UtmRJDCnoZHHyI/j+o93Bkc5y1HSTD9FV6oyJjxXD0kGSlCc7vCkdJF16q7M5xCifk4E0P731ZWB
AjVPPY9A0XkcYSovf1VgAi+V9LObrFT1VVwwTuLQ1IX7pBcPxcpkHy0EtkGQ5PcqXQL/l0yFBEzb
ZmKY9AvKXnU1nkUqQL0hZG9alfQR/FIjMuGsVmdx2PQIeRr7xlhKCpqwx2xBagdwaD6SXgnJuSQC
GhismsC/R2b/QznOrdlrq7g5oqVyqguGUbbI4uHjPIkKGJflP6AAFs6V8YHQBdYKi4neLYqMobvg
K7NBWX3TH4ZIl/w8zb0DZD0sQzvwvh2t0NJ2h9vUdm4RCL25+OCN74i0dsiUwnU90k97BWiHwhrO
klxFCNmCd+fzuQL9iuqS38jMUUNrZ6KFiga0zXmEaf833HEQYtynxiQWo8oHvJjbGM1pLG+Vkc4g
R/TeBVZWuc1s2I67W1gGw5ONF0MuvhORBIrQizC+eHlxbhFX8+Hs8gXnKw14cvKgOvLNloXiboZp
jdmXu629z0h9X3Jz/WtNqDvio4j+xX0qxa8fn6IfjHpayMpzkjeOu+zA7p3K2NpnF/E+bg1AjeeK
q8emRZH65Vy/1hZfKNCsMn5OJPymT2qwDGDigpWLfMGwObGhh41MxPaFmKMiOn8UPM9LylFmAu/B
u2cqTpdVTwt+82NNqm9HEYVRreJWPqKzrYmOn0/x6y1ysT0fx+Y2bsDDWsKdkKHyWkIdrNhv0m1B
ombWWGHrcpcq+w3OLAYgDm7BeqVxu6F3COgr6o1Q3QJK1yhG+zQ4mfGCAm3v2XBxj/lYFXsA+i/W
6ZFe3VASAWJs0GXmi2Ea7MAJ/HF1ot5E2TPPQQ/yICgm7CL+y3STJPDl7Vmjs7uLm0zo2219FdiH
0yNfsO91TEXs6H85IQUI6XI8Kqr+RmFD2aJOfWT4L2WTPlCFcKhWrisucqQslTURcmUbnNy2J8eH
PPXV7wDjvvbeqP6+4Xh3iI7vCwkAFmjNylyzEBvibNWpJhH0zPMT6Yn8fLKKLKlplRCOumxGgRZi
aXwcYvcHAJ522CrzDPquPWRJgeiq4kioE5CX/BxF7RqLHW8zHxAxAgPRO9w94M/xU+HKG+xRYNqv
JWNeQBDBYzil/qWPN53Orjmrc4HJXnJ/dMD47gdOk+WVRgrHPCnChN299YnairGSNzhUSPSHItw3
aJ2E1YpBFJDr+AxPPMScVOUwvsJf6rq2QP0iLnxSQY4WJY1skZajmerCNaf1fyNwoOg7og11NAZM
Xn0kjGLoc3vZOEb25JK3k5Ry03V0GYsNMtLB2tFh3mqMv5w2iSwjaAJZ4KLh+Q3ZfCurTZ+zHOAg
d2OXL4l9nFRcAoz5sgxqa7Osc/ywd6c2YS6pPJyCm53an/mPOrrwhkT6oiNtsTlxAH2KTQke7AdD
hRmSX2FpHmAs9YZtOwG+8jAGLtCWOWpidGFFuyGBpklL75R48vU9R9d02fDZJNkn1MlohlJUZ2Lg
1aN40914qV66qsDeNo6OM0lV1eSlSxQouUhq7P1xoBor1JKClY9JfJYo/qY7Q1u49ITL211n1ZAp
Mz0tE5DWNAGiFRM/khHM17JqZSgvCrYR7GZmYp7hv5XNqstYV2ORv5ZWuaJlzMp2A0XaRQc0b3+J
PxVTW/AQGQfzx4BjuCnpYRFCfoSe+oKqfrTe5TI+E4nQnxgCRGHKJ82RlAxdQxvr14BpNxXpAf4H
uhnIf38Qh+tWqK/b6s4h55vLBNjtcWAilj9pNR9rNHZcyuxP0nvTM+vVRBC2LPXkc+RagC7UkA2X
J257XSUxLBYYFXcc4CGAwOK/UA+cJUt7D9Dy+7EvBo/Ul5+xFnMa9tNn6ygv2LRjdMjQkQu9j5RZ
byu3sNCGt3YHwLHlma2FEAgC8BDy+VNE3h5mj6zhp/e7xqMPdM4eC6Kq8EyHAlw2HGJL9t3C/YsM
/uJ+6OQYomyDBmWjzv+VfaLlIwn3l4toYH1/qHVumv38SGkzzHyYHNhOBMajGjufVqivc2aKQAN8
IvvpZDIrNEgWY/8ClQ5S/kujw4wmUXLzNPT3fWs+0+/BgitcrrqcI80crJ4w+nm02COfAEAbIhHX
oYn6d5Z7Py9/BbC2J/iWkOa70NVEFTcH4wzpNb8Z7pL/DTQJMave4GBzaJgYKK03DPUDhibOgT4+
NCgZjqYkvWHMz88N8rB2eGqElskKHXHbGn2OBAaXu9JlGRuiJcjOPp0rGZqrhOghTCeX+5vXHOHo
lNisjaLCtVfy+3EW4HwOn6wsIQNM6FmN5JnSkWc16RkW20kPOuQ9BR1JI6wbwe+QTtRiF2vjka0k
tLzDRKt8GVecEplYI5Gc1OjmS4/X98reGKFx1SuDkNB/zA5dUGGEH6i+Csbh1HO57tSNhPRIXm78
xVDRcydkXvFDkshTRLLlsR1e7+TpsN+7jn6eMmmLRFWFcBRonb+5d5Udc5A4rn71NLWPE/EuaR7V
E8TZWAuCm335p/UTuCw0UtqjM2oaJ7NPkNDVWlDqKWW+PbD64hPNAoqeuOSZflebg7P5U3l+dLw9
QRILW6dNnzLg8S/hCseK3CL3RLcnARhVgZnqew+PjxRuU1HzJ5fuVv7AlCiL9vnydDDP6M/HuziM
xAGQaXXTPq3YTVjQfY8v714GVdRGTS2tuF4mED9H1t4qBjAueuh7iy6kSkP6xDlCiMRIw1vemW6P
yPL1lKmiG+X3YDsDbFMCKXtG5UEnhBqRwJRIkAI/Yy0HHrobNE6Kw+IZFs5aXM4CY3yIcp1w5gq5
+VeJjcCfNpxB0F58+1rSacfJA9YvCB8JwMvms+QNhR7//B8d7n451qbHGyCZjHIJjnfoULD6D1ha
9sJRVazA6Fx6rzeASsqbldGn+kBpShe8yEnbmL2lmIQ17/vTACDMGZ6o/bOVrhd0G7Yf4MzG/UWu
NHZo/W0J/DIiQdo/TQvVDoYBBuMpOdwtgreP1Uo6+qISjXyowV3EeIzSKlTgPxbjx6JLBAQVp9Xs
2QJ8XP7gjEh3TJL949pE5QtJndpvPXvNxHlb9omkmxgnCQ1Ig3c+N1pjHAFD+kTY4+G9gW+6DGVG
GPki2v/2pP1ITzCrrIwe5SJurYTq+hiVm71yadyK/alWy+EhlpwlKuGl4Y4CdnHYnj5c2BTRKSxP
Oy2lmDsiFTWwBBkUWYfoTK2zKtR+MeE1pqPrJMR1B1XgHFvV8b/widiIghopaGSqYFfcG84gZx7u
ZavfEyjliCOuSno4f6RKu3N3psPQFshXT84MZjCLBKz1B7K0kjXLpfvzE3p7w6lvSUkhtVHMBA4W
hOlhroyOtS+cBJr0BpUa9t69/K9eXa8rUkldOAVMzJNUPwGnB53nj0aY6IbSQXvXdAy6YeXOnsKR
hI9kBoGG6Yb53AO+UlDriYQaUs1QUOEVc+WgwrevlA2hP2rvTjBczaGwCctIYr3GaUr5rCPFyQiA
oLB46Xkuz2JduBLl6HbcPu0kRnxfn+7kkqF8cArQcTRbCSoSTi725zyFChEphIP95Jp7nkhjO9Tt
TX1WkU08LvYLhAhrqHCShq6cMYb6zpWEcajoeWv1O5197Uff1mf002wxtTjMTV1afxVYPwKpsWFi
tvAXHNhNhiM568pl6ZGbyMl0x0YPxg55kXOG0z7anudLy42ycM7LkxxXodwl8w+O34Xv+d5XnyY7
nI4t7keXVFE4O5LKR/YRuJ6pQiTk4UXhAhLmvhVjH6u1lqnQ8+1TqjudHTuvVOaOQ+bZL85qQcSl
KKQ3dAKLWAaJZap4bTbR/ExkfvJw54LyfG9ejwNPq0fjV4cFI+0S6Zs1rAq/XdHhZj8Eh9Gu/nCK
spSX1985vsO6BVyK7X9kKZvjX5fNGkl+s1xk6XtUt0mavEhGaGE4L51/q/ddkNthPLpMjM7J19Gc
Y3V5a8LaSLOxrKt6T3TeIMbB1yr6p5guEWasclP+w5V7AhqlzpbNmHB8HMBS78qXJWAZn5nyIgw+
4buVBBFsw1JABEoNvx8YeucTovBJdG7m8CIpG5GsDafs5rnCrG/qnARHyT4v0DgIpN4dED93vOqm
4R1eUB1dRRDESMaHzRiquamYH/tMHR1awCPWbUAFJzqN0fj+0e6QyEWxYCaptc1706cN20UzWa0M
9jQ4CyAMYgGxNa9t1wEngTeth61y5pkGqyo3UpWyBx6Gtrx98YekBItWRTaTROHtInw6s3XsdQVI
ReqDxECnbWrXqY8uZiUnUZoYmkyj1LtDMx/dNgl5tSi4gBM9RSqTiP2hVne5zCvA2E55jXsl/v3Z
KgfUCoAz5OOVByaWLVe0Mj4f6shJyBHJvQL9huZKLVQH1TiH6GXRcqScqmfpTKh5qK26Ge9IYNsK
nCoQsI9BKinmUGn4Xzemm+03irrUaNUOr+fHv9Iwau4SXlRAxMdNzX14O1jY1sq78tXADYF27U8k
YN6S0X9b0INnQWzCP2xWn/UHHqsdI4ZZmetDHi6rBMKEx2WmUqrTcP0CnKYE8uVaE4CVrv7hNDyg
0mpizwYJaEm4Lyd9ji0v/B25caUKejVMIqrbv/gVUBgfggsovNM7jdLgpdg4AaIFbFvqU35EQjxM
d5T1c6JipM23Z53cg5arK25EQadWw+2RPckm2kWXNvZV+12w7+1IuIv3uaZGGxxGN6mxJWxyLfn+
ezEtZz7v6mcw6eE4EbtVv1C7yLBwKL7p82BbebUScjH6Qyv9RtJzSm02waYbHS+2P2EPmD6z13xO
6pP+OPkkxVH9xF3b3fRkjQlHjsU9SuDlB1uLLgqvcg02Z66CipJ7jUGkaNpswmOyl3By54d8mgat
RFCSG1oaeJmpSpvJUaVeIYXSwxodB5zvI0Nh6twzx7fqog+Lie6a38GvklWDCcJ4r+An0eydIIs7
aSCLWlfallon3S5IVTQM/n7+GweXye+Mswr3ZKLkFo3qjjCTdK/5Eoe3okloFgdnk6QUK6IT1po2
1jOBif/Iku/ejN7CzsUjVW738HoGV+HLQ/alWrweKh60uNrdSQB8r7Bm8HO5Lk5MJnajW2kNAgLU
r5Fu/7aX3kooEBas54SjHv3+hoW7NrneHlYSgK3kxSISoULDcK/m6qT+3orBHjV4+VddtE27+Wg5
UsvpmgqVif2n8JC+z1hgQTOw6fH/Oy4uv6khuFs5ujt+oXKnUnargvLSZho1SbY1amA/Tymz+WuX
JWluwiBArNd8MzXpdmME3S3/rQmZm1/c4Ys+TTT44PEIPAikGvdHkHSJU6F/InFrZ1UXTqOAR7qD
NLaWaVB4nojiGXoEMd9Mx4gCCND+F2/UAj9znUBNumx3Asb9JKFIudg1bDnJTTGjozeLzPBud++X
HVxpuJ3CtWPOgAzY48FM4+F6AY8+aEcHQD7OX7pQ4JW/r725Pq1SiZMT/RV9Y+smS0XZ2TCazlqD
h0d3wxuuMIDqgpB9GZzeAaRalUyuxo2Jthbpmz/AtU0kYR2ZZIw9b4zw3D4wfTWnURh4rKlGQSzW
QCbUgpwPfBFNjxTKEeKAUE3+8yUUiOyjqN//OMPscvsGORxndKFV3UFWZYfk7iQOhf2eTTb85IcM
h4wEN3wejSyQ51UHDMgHWZ5JoNwAiXjZwEUovXQoa83SihEqnhOkp0A03UUGaciCwNibVcm2mXb3
5K94AWgvijX0Q/O5PVaS2AOCHGtGbtb6fXkZLQ3kgFRGWRHoeoUmstIdr604J9lypwZMj+gaVNPe
RLVwOZGG/aeKzkAp+7WHY1nqGaA6luguW0Rlm6MWFuNcBifY3dn6bq6xcODo29kNFFmeN4mkwwTK
lbeA53GRaa/7C+VNCVMKZmg0Mdm3BCvx2wCNpsDNP1Bluogjmv0vdOGiZgkY587IGfLDBzkevOip
QEhXfDvTWDhYPWWNFOeGUibb2Y7Ng+HdfYrKFi+Ljl+QP1r4/lkeSVa6Jv/4GXXSIpJy6uoZSaK+
cIX0LkCN+edNPfrSrTakVL9TkpS3/GKUkQtFSoBI+R9M9p6Vxh+ulSwUq4NiQGPy0D7v2bBjwWTE
zNsaG2fmcRBWoN7tf5WD8EBC+1slwkmQKs+aWDMg9fnHsndbXu4xtMidmf946g0xGppEzbY4lTnV
cjbQK1ck8KeJGvfYxFZFtcNZgC8oqAAYxMff0A72cWQzf4//++JNCdOsr9ox3OhtqTsmmYzpv9uI
8wV6/99C0SLmkhNvGdpeC5WoZVQONN470H5FVkbIBSyntuEqxFCpbtpkKYB1hQCsY9wq51fxIuJC
aEMfmL/vctrqyGX7DwYkUwnhLOaNTNAaLsjp+kisYvk3a0uWeG/76wjhLjryEBxtuW014e+ZVeKP
t2fviJCyo+q7f7z8nI7p44DdFL/qfi4YpcWqLDudJK+eVB3IabjktgslKgc1Bv8ackQBIiaVM6HH
EVseTBboQyKBzbk6avXZYkXTHJelxcD+uF9NUfkYK6I7CneqtwkZ1hat+f2ifuK6zjluJafPHEZw
8E13qvf2Bdo0RYFgKV05uTl3kaOsN3jmg3iovGCbrRds1KN6UIK58UKyLTqvuuYWCj5AnejlXJFr
9dDn2LfJVvrONAiWXWpueyJncPTxSCOt4NJ29UvseOC6OGNU37ulCBWW1GQpCX1+R0QmXsp9JskX
m22L6srzWiu77r06a6PxVsglpgA/TqUO3Yg6jR+FEpAoiVOqK5Kbe9LIiCNj667rB5zl3SdzBenf
xUqyX3EUMiiohYcft0R80Xv/OxX/QUMVwuwuvtaFUQ2GJHJMWyXWu+QBQBAd+V9jLMh/H05xHdgW
Cm9D2b9eXrhVNUjSbIKodiOyDLWD06ZkHBzTkYu44W7uxDvM7qDep4tCuoqXGk/LZf5aItAYLK4P
cXdI2fy9MCvxR19qv9qNkziY3l88slhguo/aljoxYwFJ+nT9X8HQhBl5hwegOWoq/LNlidSjc7Q4
agQ3Kavel5T+iGqhDxv3PaTO0+qQVOJQ5xsbKRUVP424+Ki+aeeaE6lLppFB85Av9bz74BAW/Q7t
EWbjvaGJO2JE9nGHsUiJl5IL4RMqVHg8kB7W/ACZSgQxwdL8vdDKMUqMzqqW09JlkTCzLa3X81/b
hd0U37fN4l44UpHEIgW5xTORaxzKevZ+FX8tZjzAF7Lz3yUIj3I5oL1ac9Jl7jlMdnDJI09ssB9Q
AzWFvrKAbJJkYh6UezrIBV6i4i2bn0f1YRWy0w7Ka878sPEL6vQkt/8Xd24xe9+R/1dizJ1svdoH
FgYEyJaUXG1kGy7FZijuivimhkWLN3++MPoaRdOSDJWnHj7BOPvic1LIPMuULK8TQXojP4mi6Pya
X2ovJa8tXnZU75Tv2RXNFKdPW135lp5EYh0bouNTFYiuAfUj3ziT9Nj9V3v6Mdzru4WfXnQunPJs
fBsrc5gHEcMbTN+t6BaCQP/nJW2c2zFz/aeW33T5iLGb0lZ2+r5j+jg72D+yTuc9rBaCBZjgHfQP
E2df7C/CMiGvPZSSNpohCzoA/iIO12z5p5AVrpG1pNSuiUYddmtJZ8FWbbVaYauztpGihkLkwE0b
SFlgdz1HhcGuG5MA5MVx1YR78YvnKO9MV1OxKIRsm+heOvpVCFeDR3lIkdOnWlOo03QUGNBh6rsi
vraqFOQMmV16a0hmgg7AShWGBtN6aXQ3yvdU1rpgKgrTJzWWQRly5WYvu6MMM3R+Tasgi/Bs/pfY
c0z2XXfUukgqmo5D4lQwvqylFG7QgPCxiEaITcg31+/9UkfreKodI+WnIPeYBGm4Ec1F7gu/FJLT
eKn7HK9t3faTkn4zmrg+rYLsw+4PHsfiREmwrCiFHrpEwfQyfox2Twtoq9u/mEHWCA18hHFIaT7N
YoCi2J849jvcC6rjRGY7JHM2v+7anOJeFbMZTuDT3SV0vk8J095c4copsbhtj+dZ2RO9C/MXX/EU
fHd8BKML5N6bWyGnGxnu76/f4w9Sl1v/GT4ByrL4iLaLqF5ISwy2OZ0284Yh7cl/HOsUnVkSVYwf
DuhNiEeLK75FbYtHosMgsJw7Y1XWNe7kwmT/2omPedGSLCpL+mjNz3yMOiDqtXXTp35VyfeRTteM
q8IHLk+DwjP0V7l7TJuPAWBJlOLZ8xt6eFLvwoB9B8d/bcj7aGdEY1vjkbo6fhxol+JDRFtHhW12
r6sq7qTGrWEodJS+iHAkopQmVll46uBC2f1XRbwbSzpdb4WD/GbwGV7mMQrrTn0JIOE3OdZpKQGw
aXtYXX8CKLLdg1f5UB4vGbEtmil5O13Gz6eoimh0hfFDYpb2Ye6mlBtLRznt/FfOPxt6PqYrure8
VhFa2NWzDwO12TkKx1TAtgg6kdpwF8IMUXwUknmDRirM3Tk+EAL5KIAtHwqj6K0WfaYaF4L9xhOm
d1FXF4iuRW9TNP7zQuKE0/904IpzwxpZCaTZVsFxmVDWZWI84saINKoi35WHsM/4TKigiSvvpuhN
RycRrOhKm/gN3BMltsQKJEeDAlR53s1RgLaJcNxr6wHbQBB9kPbpwXnVI/9ObkNwV2RzouduscJo
t91SfUYa9KpiKNarATVgV0aIElF4y3t+a71HAJNZV2lLuOaMcJy50gfueaTxWH1zSZzI5y3Q6IwK
Gcxg5xydKUZE5l4VZjId/1YLeN42z/+4xCFgJkC3R+s7hvq/kDV4uxHA/GoHYFvrtprjE4Dt3UBy
ChE4MDMavaI1sh4RwfxtlFF+lJFdYLU27P942ODUOe1hydZ9Z60J9FM0X04wrd4C3ZSVYIlmYokJ
/oEqApHS/tvqrxRXFeUEZoT3NO/clk2B7C/PWPck+0O/D8fLSKehcIHuiyDTAIyEH6ZTKmuoKvMO
pw72W8D3VtoXCwX7C4qAyVmR6H+kWmtnmHKGE2DoNz2cemf6jNMxlmPsCNH2Al4lqMglicTZS47e
L4uP2Pl6A5SxcejXP7gkv6xeCk0PHBQtR/2oEWY3A60QNiDqUZsjFE3/0mo6JrABOZfKQ5mXAKes
koH6FoSIY15I6HvBMEvkDQfQbVDp92cDydH/cQ79zDs60zanb70ruArd8mBxg5FgKEhjRRTBwSa5
BtGwzrJ+LTSyyFBbFL6NvcXcRTU4MHKj19juckegp0sjSzMQqST6B+XK0vGP7EcXsW45JuICKYOv
qVfQHQ48KEsgzmECum/IEhSFLFwjaSv4Kq0NOFBppWNQTN/ZcHfVZeBSLxppz2nGEv3Mte3IUTCw
SG9V4Cv15+sSATr1HgZbzB239mbfUyqCki+qWmfvEFtP6ib6jAlzXrtwbfCR+omThMyQqtLef/0o
u4C0fV4NYLQQdy9IyjP1EzYx4qal1hAB9toWLk2BwQyg4v1QBuFxYiqow4JaluhIo7/K9djyBNDs
2gmsnp1XUlThSQcc2k2BmEebPiCRzr54Ve9znAxAQWkji7dGLii6EXafvSe+jeC9FiAckrnGLtar
wdiKd+6OuPZE6HoNcK7sr9xo0VbPCN/eT5fq+J/Ahkag4+szpcXF0KMlPcA9pxXrHizRIoujXzpJ
aMgLXTt0ueOYzcmX3cnDtl/Lsa3fAvxn9zb3XoQrlpRCcgBWnb0h7oMsVkuLmCq5fh9Prr7NlMGv
mivIBsoMwavJ5qnfttixjrGaMrp82ch2QEoA2pvv0UYFYlvD9GIjWWz+r+x1LA/cNuVoHe6BMQNm
L8XOYsPzpiSCB3y6dw7GguqVEX+zDIdy3+LLYLjCrTT6LKH9QRM1IG4xDS7aIEGUI++6Cs23fpwA
wvgdW8Qv7LMgcSRjCtWU4w/gSgmUO2boNDcac9D+OSXzeJD/6XPLZEIyetOWwlxEHoX07LoxU9+B
D+7FDTiY3EubRlf+g5/lvAgV6pb4nxlik2Ei96C4rQ4teIfIrJCopnVghd9ogppx57+bTUiA9mZA
SdhZMUyZIf2lDVXVWhkw8ofG7dgt26GPOXu3XBzIhvG4Wlh4trp4FZyJR1G/p7GAt1UpOOc3D777
KQZdLcXgWLz+yvHxkNKjpCcAOq1rrW3wf22WZY+uqhdB+VxDYz9WNGtL8nWfCM/SUXHhzRt3lcCN
fQjz7cxvMWw8pDWg1mBRb1RiKrCxVJrPaqc1phfEiMsTkC0sVexWCAMs9R6Q+AUxqp1BqWrFKLpq
3l6qjUtlfFMlYdkJ64j1ykUFbSWLUQEpvycqtAWDTuvqrHEVfRb0mSh/0Zg93ngLYtN8Gpy0XryY
WauuCORO5ruo/13v9AXMMMDPVoJla0KYkFmwZpPlEkXEzwCAUuCv4A4NxP5IFHmtjuAY0d560RJ8
xFouxrLDtkbDzYdR09krPFE1+hQ5UEXP2r6DIA2XCwwWi9fpmDf0/RvVRuOA5nMGzuHyVegntNQv
onYywlAi8677uhsgWgGk47JeBaeGbU36lhkDicpcVvwUAPNvVn7ICrHzHGVtNuTuP+FfilmlHu8M
RDg6UZqpb2DFD/KjOegH+/0r+ABxyrb8Soidxwh5HMTdP+mALmNdQ82SygxF7XV57j8SaHySrQqe
Dw7SvsxtJALqEmPke18YNcHvmNfNhvAVVtfX34ySU8AgjEneso0j1ZyrLGlldvH2vndT3dpjPnA1
trYk+G7YbaJPz7GAYLiQ/CGHpKOXo3BI3Dpuw8HHJVKYodd7EkWwYZLkBHTaAw1Eb/NHwiUoK5ji
lPhjsJ4Y6JWJ6KeBnc1CuVeJTaJvC/K7zbtwMkEwzGUxHel0RACznc0aBimRpjzVWkd2zAyORehy
KKowwcRD7VLHQS0RFRZAkvJK0FVG6XqyhiYSCsNlbGsLxk0UbVvNY02VlqC7j3NHJ1MmOQkaZyP2
6lAAAXuOrp11jp6jkJqmO7z525OLJnpplIKMcy2T631Tek5vROpnibrjb5jAAy488cuEeKGL50ds
0LtUIQLCqP3Te33fEIoW72Rw/N7EeMFVFlla3aUIY0xa2nfb/hwjWHAKRW1t7SQNvv1j1se8T5yz
ZVPRSgopIB3dGQy3qIgYdbSVEKXuyJP6EFEW5T1mohQ2LpoFzoDOvSuyKE1bqpBQtdEY3bIaw7wD
avQyRHUVZX739KTCnAqTlacNNhEDnfd7/LTLQbFtquDHTrs3C34g7o3jHReixw9ja4pYESaYXYy4
ObeudLUxD/Z/8TJxUE9Dn0DuoAmfFjBTO1fK1d29ogU76rHxtfZXkJOWbjsu0qDQkkrNSxSJzDcU
XtqXwuNkqVzOLwWUqvrJGddbKwbhJje8stXNwfa80b92F3bJeMhDCngmYI5wPBryFuBz/vXMV7vN
nzm6KN7YkkTbBvs1JjqkJHC2au+gpOxBQ+YoolwpX87GMvB77VOS+8PSHCDN5HTO/aJX64nZGmgT
EBeP+pveM306fJaIuqx1Ocri0Ry6h5C+8Sycen9TseuythmZuhdVMPvomi9hxkqC36OJKzMMFlyA
SXpwrt0l7FnWJ5SDeXCFpl8G9tdErLdhV9IR0oe8RZZBJWr9WTsUWP3swqF5ydK7rearDEV6bhK5
jwkiUBfzn9bxCI/6+2xHvWojnGLsHbsH+rS3m2ug92osSgFwmUEOk1mMvAxL4go4RzpPfA66CV1o
uF8Tr6nF0WMPuzoUtFKcgaoPodDJAA9nAOju3rrueiwJh4meFaYHVZ6rTLiaa/e3wIbU4vMmNfP/
f3gSLsNXx1kUWRK5hK+a7MWzVMfb3JD+T0S5hVgZZ1speac2UBG/lJg8x6EulLLoxZUzPkNLvSru
YZ5cCiQ5J5EmtCPPU2+NcH4s7qwmLEO+Q/C3+orPtOxQIcXNE5jVGjqegxEEnB6oJ1xTbw8MVfij
nK3HY1ARYgEzy+cb6LOEMM7ag7BkSbfdgl/+uwlLnxUYHnuLcXfbAZWLxX9SuSrh50SB9eGo7+C3
VkRn5JfkcDq+CrZkMWRM/iP+zezq14DERZM/5Rk7e4lR89Xv7JbfF/DZNCOcmH6P5w1cVztHLSDD
OuQ8NwE0MpV9yo0wFSvbZ3HyTHJGEa0Gnc07MlNsaG+4jg3ZM1HqCDYTvMm3djxZQYxNjRNjsx2J
BnGfGxE1+5fzItZvwUIT/zG5hEtvX8alI1jSUB996ZlKmmCmN0JofMZL/hSTIllgtLN4RRScwb7F
XHXsyF16GcBB9GlgYFun+VgndyYdbpjDB/AttQG6nqh4ioT7EjYf/dvWdaIitUznw48VE3iSsQeP
doQto8n3+WOCIWWk3JxqstGaTse9FZjuxjLuasCFARvZ6fSSK81OhZEZc85q3xpqTuO6HRYNPIBx
z4eB7N0zwylMjP3OUZuSjRM4kpETiu9kU5g4Mou5UcjNgZYlMp0s7oIzy7M9ChnBqUgO4pleJsp9
xL7HBILW5xgUhxZA/Y2Hck+B5gDFP/fCKp+OrIUaO2zoK8v8zujraJs0w5+3ceij1YKsGdIMqsdI
BaYv+2iHI7DA4NRKhFF1I8eZxKSYwv6Uc27gSWTeeQ5nYczYdtFZ4I0hb1GRbIAKuc2+ugK3rCPy
0p6ujH4Wj0QkoYMrDlk154VM2D0anBpaGbXFjfVw7gdSm+Z/srUXdnHr4JQhohqL51ea2+O9mtyQ
oRKlasgeYAlvnvdtx11Lcb5sD5A8zKMLNO3zwGJ+yMjHXBEltOPknDfGM8SuRkbbBRpYUq1EiqUz
HKdNQRGJYSeG7qU+skCglmNDa2wLnlddskCw4+PhGM4B4aKCNXS746u3WmNG1ozU6VtEGIU+IxuN
y2dN4a5pbxtHZ+xEpIUGQPocGvckANpafZaD5t3ne/ZeKT5mSxB+dRNJ+rL7ayu7ozUmpdFHsbh6
+8q3E/Xth/4/RYla1D0hgEpOtdkY4Q1GrZ0SEQ0LhXkSpbUN+tYfqEMowSHsHO5E7pCEL5y83B7v
mmlWqUp6jX1F1nOQF+DLnzjCrE+glxiGTOd8TMGYdmN/Zec5B0OkYrUjEruHu+yPtQB+SbNwbV8l
3Soi4Bz0SkQjgLI+fgn+psQ49zXub5uRa80eRED/Z/qkPMrrW91W565D1I0E8VeOiJ1EVmzYWzQG
9dPjdk9v6OLq7r0GCLHQRSqHbtuDe3SCfvm4B2m8VoXiAssNhxxugfxCgRwGX3KWXwahY4i9Z14+
Otciu+XFHeH5y0/AQMHZ1KlSIvH0T9LolQAO+VZtK6RGOZaV+jm2ircP6AAxMW+7XA5LNU8uBm0x
Kd9FN56p6/qrUI5MvH5tBku11s0CX3x3iKeqCPuLPCi4a3nVXLaOaRP0OtjTvxw1AHIU6ObDRSCt
EhIYEI2o8XMbjanbZIFrpIgA5yPsUhXWC3o5SXFk9Gj5KnPbtBlPCWIT/RPU3ZUFsAKaVVBkQP6G
5UheJH6ySuE9NWnpOZktUs832oh9WZtoFqRZ26+6Nvm7+Z9HNJEnoS6AAP9g8tURDbksGn60l/P5
DztjGmu5xOxfusTzCmiWOQs2lj0oyzyWduxalvD9D54nNGg2XfGT6bNyjPBqqRnJ4LCb1NeQuXuw
tE7M+dJxE2hKLOSW58OHz+0j3cyf5w2rDpa5OYYN6ji5MH4jDYVJi7v6y+j3SVaCId6YI34a08wI
YPu5P8rrDqMrGE71+GuKdBrAXTl7qi5A2Ny/DYVyR2RzeUrXGlPAwbYZg0psBv+wDU9uZRNI3VHf
I7GzG5yZwQCLuk9aLf31vG10EU8x2ZaXoQp/pyLe8vSOPd1JgeCxvMZrt4OdBjkx3GyIuguvpwTQ
Prsnmt+bFF2XlWe/wVE/1Tp/JWdMv1AIrrNjWbnUKGmbmT0oZe9AgC9A7yCSP4J6oDFhVxlWCzoF
R0Op4dDQ4cv0y/TGLXtL7nedc5ugbqWF416rMIw/nI5ijCj6lPlrRZEOr6qRXhlwqLqYohXeyBpP
EX0d6uG1KNi/lG2sWGHI9vqarcdHA67uvPpeWLr6ZUlBh4UQ/g5B+Zfhkdl+Fqk9XNApTobSh8b2
f5nO/JQ01DWCRjEw9hcc8Tffq4YS+rn8+k59KR5p/ggd8Z+QevbZq1eyKY9A1NEySICDPtm5C5DG
EeZaLan19fInSQm4mgpeoFvarqbS0rRFrfUEQ6t0fk7HfwvzVeSauGyoDTRBhXg6hqcOkKtIyVCv
Nja1Gm72FJQ677tiJWVfhl1iAs9qTsZA0JFkzuJl3n171oZ6HeglSepWE+Dgf4cjb2yObO/ZkviO
n1evVuZT6zZrKp1sN5Lc+hNuhpbjDi629+TnyxikO1kW4iQAMm3M86ROkCv/LhjCfMPxuHAM+YZg
GW/kfj92c0Rv5MFZ3dmO62jTeYrcaKTvVyI5ZeBbr0WABXxMW78p429MlPr9zRH4RYl4SjvM9M2v
OoKE2sC9sDQA0BteTl1SsKu+11i83A1cVW5ogNMMewGbCn9msMQM5m0zNXR6/IfqJxXfrIz2U7jT
AHjwuPzfFA+8T0bSvUecAYBMdU1+z2o7ZgAgBDqz432hbpozBHvrVFBHUujMXGRE81qBpUT5xJyv
Y5YUoMMUsitjvqi1cHA9F/0nxVWLNu8fgf524/4MQJE+3fCSydb2DPFZ0DV0KF6s+iVfnzIkWeRm
7U9HIrClyJNfHvLDmRz8z9dx9XBHbIz3yXb7ij8OIbL3KFHgnIxVkxBmfsh/DuedmEOcAu5h+K/l
sNB8MYSdeD/FNf9M/3KEInExOglOEE3EYY8WR6r+d2/8ZG3me3Z8JJF5MzTssOlrAyrcbiKHVe/H
B3Nw3Nefxo+plSTaHqGH6bLQUeX6CGqeiLVtold1Wn/SD6GmVMKy6y8nMt0Qt7GhWO+Y7dQtphid
fj2CHjkAUGL55Il99A1AtbquTax9yaXDf26fgz5T/ksCcXuYaOmGT/VZySyg+3TQ/bBxkWuKy+hi
Hp1FzoNmFNn+JmPqnfAbKWCo8gf4LicwNPwmmzIjy+1R2NsoVXhP2O9k7Rv418vBRpEZKd29ts+Z
VUGhSGoxaRm/O1GbC4p54jUDk7kYFpCkj1NYG66T4Zvf6vk+8iuvnYiQ2D9x+WPj/IvJRUb3omCc
vf9la9KUPODZT1P1R6/0yBrLRAwh4K0G/+5dmAp+AptRrqmm91SbNZ8Gr7pSBnRfG2J2OeJoHKbq
/+WuVPRFaupOQ91amH1YscGHBRsV0kiz0SRto8eIiSjoNFTpx5zvhFvxV3KqExiIYKks/Ump3HWF
apu48K+ZNZuxahVCv2HZRg5noIKQxaI2JSzGmvJrr8MuWZHCG2nBRmMvTFE9Py34kSN3bDnPp+zY
PKdSCsB5JuOBYIpIN2thrPDBscsw4MQ1NnNYQe4JkmcYt7O5eHWtIVTSSv/lNlRueMhVm53mmXaP
rqIZsEI5P3jk07+gu1HijeDn7pldEuaTwGVGz6B84rXIy+0vvLeoVSlTUg99aqgfdUj35uvvwF74
uyqxuGxt4499nwxVAeT0aJDuj7TmcXhhGjLy300ODqzOkYu7IyAw/rnh+rxsjTy7ddH4nVXMa/SG
M95LgyUfIzZWrcuC1aGMLkT5w+LGM/Rz+p/9E65Utth7pFU7SJ5azYVIJ7SufFPqVxiApVLrzSS5
az6loXtdZ8FQK8AqdZdmhwlHJ3iY7T23f8Rm3JBsMBI2cbu1UJyGU6iJqyIepZmjfGoPxK/nQdco
JEbodXBNtePt/p7moTYUHn/EN7ZfuNiuLHcT5dSOxsZDiZwhtIBfg1+L280+01qYNKtsGBl4KKFa
Z2zeTf69ErivZH+EPK7IQB3qXMlxfeiodgGobXXA+q5fy3Z6jeUsYKx3xxJM6IqeWgAZB7tHM2Ar
23O/27ezBqjSC1a7y14R3q/s4fZvJeKhkkYcevuKtZjr4mkyLDPNYRh1WKR2IMhvruJ6RyPUZS1a
ZXjYrUdEI9h787uePN6GcPrQrq8+QnBg0JS1s1OfQRQLFJqOGPkNZNi+67g6qJcd69w6zkfgMPo9
sgygsjXluyHE5raVcQ0DroeJtOihotCXdvTjzIs7Uz/EjdPop22/ZkrjOWT6p9wxne2TntoG3K4R
WJlMSN1tRkFDRN4gcFZs6NiBPFKP4vw2V1GpbxjQEm0s5PI0mrimHMWr8r2635OEVY5L5orJvmWg
F2P4lfMVba6Jaf45KMnsfA6Et43L7u9IYoNk76uLt5I61zMjH18eUDeo7QdUy/+hHOHQRUpU4Rkb
RMw66lMaFS25UxdQTYTZsT97RiqgtipZ5p6GPex6chd2ACsJ+qd+t8t4iYjBOZQOKfW4q52tdbGq
vuU3R4xAnCogmGd3g+DaNaHqVxWagJmzdCBVfnAdVxj8uMJC50S184WENNRq48useSImpmCHH+0j
Q7bO/a0s5qSpk77UgP2Y598QGW+ZawKLSSspJjOTjkNRk6nAPIfaqFBucl0UBijldfEGw3SWpWX4
JxigBCY9mf5GqIIlsLffdCg2B3tu9FOtZwep04bJHw9ZbxfEZeX2r7JOiGHUu53ueCk37qnAk3ze
yMT/63f66IJd+rbKMhEKft9HQN3Vv+s3mxU5G1sfo60cNwMmEuzPeVFMCuCfPqgTyWxoPl3BwEc9
zvWumu1lkRanOyvMboLyUuvRkUOIjLVSzhPNaUSLCXeGQyD0qe1UzbvHlublgQblBbbzVsBsz/zB
5K208HJQMEygRsrPVU+SNoOHjuiGLWZFzDmBaTFd3YpPuNtzhkBe/oVY67IqKZS8503q+FO6W380
xlbFYGqonmMn4U+i0OEBnJDDUfYp6jzEd36JyT8PQFgVSU6duvpmMQ8Z5d6jayRuy9A58hffDWgC
8S+OVSDH5Y1TJmXjE1lt+0WiNFekaTDRrJbr1oZQ/IbQj1oFx6sjuMaL3oIpyHvykyH9ncN3HFf3
90pPait7NmE6LgRqLW3ffG89zGcpsNFtVOKzXWpuWKNrodpY4D4ROc6hXrvWAJThIYZGmKXRe7tF
zHqYJrWF5OLezqk5yqjMmpVk8vMH6g9AzAYkGpkYQPf/pHKYEQz1DgR2QxmAfwA3TTse/l2kE6rN
v8u4eI1eFB8rVWpBR+vwptS7tCUVcnWRuvNGAiwJ6SqozCHuQ6emvZsaq9LDmNnP5OVzHV5Hdph5
pYzzXs6mtaDniYgOi9UqqsBIvG0DZFymt1HI3yqIwwj1DF4IY6lkz3Y+HymOrDj9XTPSUo+Auohr
nn/ilnjq2FvfvYMMAX5azNWlX5WaDmDmo+1kF9E3HuOxYCI7fJj3k6WIscS3kd6GPUhYREOZHVMP
qZ/lDQYpbGlOdeZVwZzgW8AaYhbUy1YiOusjrhWLWpHJq1tsm0AbLVrdUu3stLIpbACGTsSPKUgr
ulYb5CtLsrZOaRBtdCnF2KXCxmBdGpbPVyn5fx3wjAcilPFrXcJepSB1n3ZHW3NFWmcyrGOVxo78
ZRwzLbb63sApvwYR7eYmSFDeSilJxD/YXqX1P3No45WaaJm1Hu5rVFP65cUjzOX+CEwCtdnddL3K
uLH9kLsB4aYdDhO5umAlc9Sq1NFvGoy+AHDWrYv863mHD7O9nU2mC4Z8r+SslK7ATHCgGyL3Z4xV
bpBRidaNnD4c1d823Z4O0DphgVrLWWejezIr2fEargiCBvUgnvpQGy6nY4EOLdic8VuZEIrVlx97
zp6HYjRTn6LbJpLTybhpWxDP3ffL265ke0KtdTBWGuJPuy8KAbzIs29qkwvf3Aq2wLydv6HeNtsn
X4FqbCgpYX0q7kvUtJjMDvNLFrBfg4BaRSAnQbz21qGlcYd9ciM31lAcbHaypls9A3iKMgNAz0po
IcDlgIxa3+bhycJUB9oqFZrI8aJt/F5CLNNdk4UYC+V2xOwm4fw3PrEFD8UN9nADCoDRgZ2aK/LE
RPAFeNfzo8LcFSe0gJxQ1euI8XO0QbLaXL91hsZSsmUZIMPTkWWMZin5eRJHOL3MhIbEsxBNe43L
+0kvVsa02GVwuDttlocjF67eqXi7NO0k0YwS2uvVktBJd5PS0CbLID+jKkcj9W4us2nj2ePn2O7c
UfomASdf1l3DxQso3Si9M5AomDV0kFhAHaudHCnnyR8k07PLaSPbVdwT4TobPw2jZScalMd0yofO
e/3YbaI5UZDLrdxMdBoMskWuwZeirzmY+GpilDFjdWzwclWwEp9m06kXmZ1kQ19JtL9nxshfmH5M
iIhP886xc7IP85GhRyNBLHA+HUZLGs5bYTiUrXQw4ILSp3bEpl7V0eahAvQxCAV7yw/wSFbjeqRp
bVMFNh2IkcekrLxFbnnDgIIFJX2wj6ms7Sb1vXlkjys1pLwEf8C1e6nOlomLpeoX+jYdxDnXIjpv
TfoF3OYZkQmjv1ae3A2etiqvKyFypnI5GeZR6VJCVDVzzD1jTmhlgGgHVyqx79yhy3pB06UThztt
jIXIS7zipt9yWiwC2COvGFOvgjQA43uUKqf1Aebd/TnJL93RZ1qU2OMF8PukYat9FiT6M3rsK0Tx
n0sgYO/VcLvNE4MDwR51IEV5ruycMdcZ2+DIE71Ct+WlKUD51QPX79HWiCjQ+omX7tCxeVP03ZEI
TVYv/tlN6CLg2h4Zi5UdZo4NRokqdvPE7qoFlv8ZS/kkjvyePaD7dIBupJr6R4qXvxJLAGgFKh/b
l4qTxj5VytbwqJARQErkkwH1mv/PY1iCqywQ3E20/0QFRWr7Ru4SfWxQMynq7yDAmYUU0I+sfutS
Vcwv1sWouPXGuuHJ2+SZifTd9s+bKQX6sHt7+n0IOOsyUsSoLqYEWxUhOy4gsWDseKnqAPyDj+3R
qOFvHxBIfvk3e6PU8/MNhA8Qza0x4PTNfPi2z/4F24FR8UeYQDlrY4QpI0AGgjqHI3VVYT4wLVNC
mbTYGiCnNk9EQzByOo1HTeaGumvSRRUlZlMopCpll42ZE0dcVXNIcJDr8hsZcGw/O4xoZZMpkCup
2m0sm2z36ifvkj3QIssKavXhNAN+I90UoFbVIKcAfWqIlKm5YpmC60vPT1paGJXhWF3yWE0VyUAh
KoPzGuauAFCL3UHWCft/Fuj6zdN0j5EbKgWIIGkOou76LaKN2Ml7RK2RB1PfD0Xy2EKgcdxjUTDg
+GilzdEv/mBvZxyjMSGW6ltP6PoVth4mnkmOS/ajrrQEKlWE3RrA7JKOoJb4q5dEJquGChIbeZxY
zekJkwJReb+GAxMRf7foBmQo7Le/tGLdwlckR/xABPCCjwRFrILw7WaPHk5wO9ycYRP+Qgu9e2UQ
Ta0r1TN/Z2JVZ+tvo7q4fqUnmQKl55Tf2Bzm1jCSEiR3jG9s9ArUJSqJm4lZmSSUgu/DSOijAMm2
/d5fBlpryj5BAxs4HLzjz+ryXG4Q5yGO6b5da184P1UDb5Sx4cXWKmfo6BRVCiZRd6ufdF2c7J4P
fmkn5A9QsvkvWKxJrMBq5LhXHAThmcVyVEecB4XY5obdr7lqG32RbQn7uxSzH/vgrurUWPqXZyog
L8Hanl5TuK0uQ7TWbGm/7mydqqbsVGg0XO+MBPVjAkevQN3ncSmDm3mR1nXTgjPg9itOnMIKwnxK
+YyLFI96AGaO33GBnSclPhHIcU5REcABtWurttHkhozwIZUiDS7fmesmAQm48kWaC8SmcTxPl9QX
2LnnBSJj6boI6GMuYLmo1svF800CjGItyxP/xRJcQPGFqn6bPd9fg9/uteejJEC9Id9J1iUZPq+S
zTyYyZ92WwafQgKvyDVUx185BVGxGGtHWgRyQQwZ9CsYjdaNZJaN9Wnu9d1O43FJqB/N5x63qbRC
JckL8PjasgjO4GuHEYTFebHiS7593qFtmlaggoKBoVwja56NKXYjBHfew0a3kwtn6X06bp2uCcWW
XARf75yE2ijAWXe1Rl6LtxPHqALnjEiqEiJjgYsiyKo7tYjIgMT0AOQ0y8zddX1xQbjWLaNjgApK
gbN31et19/y73sl02beCwxbAyRBZLbSRvYBPwp/rqHuVLjahR7ZxRf69+iZrhtVXucGjgDfTECzn
/DZD0LIXuDgnVt1kw7r+YkMnAs+gU0NGZjlTJWCLx/YRU59WyHwWkEuj3BdR8EoLWAzqVsjiQ7aN
Et2UwDh1mWBB7+jM89DRcDjL5sKYswG2DjEMjkB+cG6hKaEyYNCD+w766c5Bx2RzxyKDsiJcHuy6
0+mij0+5tPv7700xp7cUSqhhOeEbyU+SK616uFfy43CzvGbimwctDpzRxZ0YcYfeK+sxCKHYeAYG
8eP5NgkF721kO4p/nE4IMbr7OKtdDhkdXvQDqWsTK6ACy+bvDkLgU+sSdUeSV3MnoK8kNA1ztXJp
zjTeSGAfOWVYMHtDXeSSTfHMUm9pyCz45VIF6MTno7t8GeybrJqbfGQR5aLbno1wgFuS5vx5w+Vm
RzEgRLbPo+IUMVialgqO/Q3TASpshw7ZO0ofbXtOt4mRWqhDTbtyw0uGIDjE/bxmhxfDNnn8wX22
3fXhwQPeVU2JUc7zUH6h+s1fFSjWr628sIQZEEoUNKfZh4bJ1kFJZfeMwTGodvQqi4w+Fu1QEB7c
SPSF+/mcQd+TDeYtZLm0QgC7ox0td8XrqLbmOBzniGvliKv5gaWmMrkHuRIDUbGmOAmTXNu0/Dbd
e2b1K/NxEgrfVj3/4aBNvuFZkCBp5dKLBI0yX0Al6y8pue5gpprzN+Xxl/QbB9VcnYY+qJ0av0Er
A/7Ua1NO59mYcRcKeoZsxgfzuSvtioVeYrrk4OlfmojZ7hNZ8wE8kx/eQpt0CHHxZD9vlVOn30qS
Q4eopAUAtf1W2K4xSMTfHeAeJLF5/ka0nfMCAJpReaH9HD2EQXlmuJJpO/Qkp3Ih4RMvdjTpZ7Z5
7XxZzGksJVmwiPnkWjtOZ20u7uc9BDPVCp4aSLAqm4BOYBNMMoxolMHcKbQOH01lJYwRm1DFF/HQ
6vurTuPPNtsrBgz73m1iK1bzwDfKmlv4KgVBLgf04TrFzTV1xFdKqaz8KsTnFXzYmJ3ctlENUD4b
D7IDQ9igxewspv4DDqSaeKyaAcVD0pGnEO6yRo+sq7XDMfx/WPN/lNExANaSXMDmYinoIQHmZK4H
0eR3GrMqK0m/is9hfm/8Lm1782xhGX2WzSV2wwftSnA2jU8BXCv2/X5aTXN6/ZyuDHrHgnEy7Xq/
k8LOtPgQ0Nfu37MpIhhBejCD/kISseFq/Axxn/khBilvbQBwdu3vKQghL6r71i9nEtnoJkcxLEyS
dfbAtSotJa4ze6JeY07UqzTnKeQRirRFLDGmeQAiL/p82idxTjK/bcNKd8Gi7oPxlUqmxfQ2rifO
TQ27DyET7u6OYsbvwFVi6nbFwAMAZELZo8kQwjBDJbx/42CtoYbIuD6GC70TjfxUMMbZb0SvwMY5
I6E8cHPFtvKfKVeCS7cb2yeFJ6czbxTB+jQ5CSZxmS+dqH4nRpZu7Smam61566DdDzE1JNKnPuq0
sFg89hx/78+rTj5evI5EbYiNihvzyWv5NEN/p77XuaUFM0AMiWui3vUINEEBMWTm2H+Wjo9mxaCI
Ot7Y22NLtPRIHOLlBbCU6ohdYcjakYOXKKDV/LbdLcwvD+zP9YWjIbAJXqMZQjRzRWkinGh+KLcG
Ym+IIt+71on3Tq6VPq494lYN8R0EXz/NQCZAjCqCpTPBL0vP5kxpDyJdzqHAFb+uwUHyTTmXLVU5
TgfJ9Pf1m9Dx5V1NlpFjBDm8y8VA17zGe/7LaDZjYqkM2sAiTeOoyRlkIePWpF39cR1VKvlZyvFy
/giJ+2KwwG4rYY4DBCRnjoyOYeq847oyWX9qhsK+is4V7mq8OF9JCWb6Rkas0rg/+jQr0zON1RdS
7DAhZ/Y1eRyivji5Nf2HzS80/DvFBWg/Hb2R5apnN5Ug8b64GFgITmProp9GZEprGzb+QOmUF0j2
y8ZOj8xl1QHKk+zMgfd0L7IphEMALPz6xR/7JJHf1kEcae2exOgPpI0xG4TwdPCW6vQNXCtQKeTc
ORgvXaKK4YxRDyogoesErxp6uurIyT6ztodnKgGs5Q96A/8FJCTTD0j+/Q5vVxRW2ElXyMoBHuXg
Qz7gc6WODJ1nPv/XME38EIgwG7FIr+zab4o+CXCqyguhY8pBDz28IGNSkKjThsqV2cgnBp9JHFQ0
3cBJp4ZfrA94dyJS6nNGneLMH+L4fCTU2bI6EPCtK8rJqMoPMQrAw5f7WNjDESzyazu1IYKR6e8L
G+4gsz7RmCzDWQSW6+9BMCjhHO3vF4/x1HpFcIx55D11ZrJWhYfltdU7W/cy++GAf65tZILy2jZw
bWSmt50u9ySSdVa7KOJaNxPyiaSv6lba56LZduT9FroULqN7idsJskROfFiN331YUVx8kSPaM+SF
A1aHNh1MhidCWZACisLqDCzZ0x72JkjnHnJazU4twrsBAiEWCAzA67jZ52IyLI34W8GkdIWuT/iN
p2XpU69C6hmiPF/apFKb8jLY4yedvfk8V6NA/JgdITGsDC9hXG9aWtnWlTH8QPlP3WZL46ztdXo8
blOvmyiy3p149gvlbs3OoIE+QW9EoF9K4kqiHg7cTsScoRPvG5DonGPTCOkutv56FWhuJ3JQAZhX
XSv4LLIlvXfpzNaxSWpbzYs0RQxitFEN4kyQ6d0zfQyeNsSswI8ZKVC9u8o8tcFSH/LsaTbCcwvC
s7MwbEaZiQaGAMSd7nI1mxxIVESciWtG8K7pbAYvF2aufSZwD+01KSIJpc0W8dqrw5sAkxwB/uoj
3uH1vUHuOKp9Za3485v3izN0f8s2DWcNwN3oGTXl0BhqiVK9oOMfjoiZ3VHgP/yEgSjRhk8SM8bQ
Bv6Y0Y/9hBiANJr10KmcQsTuCOUCD4IsqsL2eFglCzr4pHYeFuLcJFSbKlEoM7kG4Hu2LGGH8SCO
iFWsgPgKjXDx4smyAWTYMND70ewBh+017qbBslx+4Ax7h6GsWUA04bMk0GOpQu/o4V5K4DkFspNO
onuyRx0EBhIWMcCGFlvG6YlKNDB/KeL+16LlmPDeamjphmBhqf5rfYX9X6jd6wjobS3vrCn+FxZ5
2LuCOyBUTwlQuzJ1D0wg4xpl/uVeU11UR5cw4uM7v+q44nPZXltFS1JTpdglt5cmN9U3rztHPmZT
BEr6XrxTTN2G1SggHHczEAua7xkJ6flN6ti7wpYnKeyGsm9PAy4WriEM8QdnfGi11CpPkvPQBdof
pA6Poirpkl0tcstLEbEEx6Ce/NdcUhGOpia4MDd2JDV0RrqauZ+CD52Rau2a6WiTPJpFSrJk00v8
q9uHQaCcD1/iixPuys8GiwRwO/fxKsvAsKoD3oRlf+Cd+MmS0qt4Gf43wNMIDYpfcgJEzDjVR6dd
EKtx9IrONee6+EqavJBG3+2Y8dTuXcVqyeegqt8se35Y7UjLajBfD0XAKRsIgnhCTJyzh9cqNGCT
G9uwWMvPt/huxd+Lrsx47AuL/qRKoIepSdt0Kqh0Z4AMdIeLaA7te8ApY9nzD/96cdzAYteCTqpg
5WPuRrb29QsViIo5ghMkAehdCbdNzSu7emf8IffrSzpji08m/Jx93V15HjCvemuJXmDEYWDX6/bs
0wdg34/GE2JiAmdmTHQl32TkwKZJ7hTDzi3d/FE924THgy0WVJQrXOf8h6VNWQsjFHM2maGfcYv8
H6SobDs0NudxTT4jJYflQiAvrGUwRHYzdY3LEl7D7wpOLy+qOhmBTs8XMaMIS8F+QwJ2ypjA4OKn
+LzoYJUrYGIxYaKiBZVrsbB119+sgN5FCH1XgEC9Cl3B7xCKLSZ2E672qmsmSkymm9OrGwH68LaK
QbEXR6zHSG8RjjuXPv7szgX9J4mPeU5Agh2/TY7MAwXjUNABCZDWfzJvkHz0gl/oUtY38E0BEjpo
U/a+ZilRbTvjoLvU++96FX7NUtk3aDw90la2KovPzwuu3H4EUqATVqpbVut+QgoWdO9sGvhljR16
VTrpA3p48CX3uLmcm7jtG2oYqb33GQuk+AlK7IJBhBouD/iDVwCxDA33dVH+zvpa2ox+3DGKf9vT
rZ99QUnWBzoRMdNwnEPSfZFjZUl5R/Uzd4TjyuYF7kt8YbKLBnAuGhwYK2agAGy673nxNN7TxVit
qlv7H+DRtHzNWFlgBoWHTjiuqM3JAiHwQsSNwt458TdF/tbr2otAgd4a6zz7hpasxNPqtogmsN5Y
jw8HnbQz5Ljf/tqt5nOFahuxgNQCo4mRFivQVh0atO5Kw08O6lj/iKZbJ5/V7RiKfp3LxlF+/g3O
2/w0agWinMd2TJdeWJMkIfQmewAvQ1kn1A4seVKReUsWInsWMLXYAZQ01sdgNQp7sWlex/2A1ZpG
CLFCVKpBCktlWrUmgl/oE61yEbA0fVRxCHEXze2ilcEVOJpGdnBjfC4YNbeqVzeVr+rD4Dl0UDZJ
hmUNO/RB/hCiJQ/d6rzHQ6mO/UNeZIFAwpnnzQ1ajHxaJ37K0hxIBPRvJU5KShDh+XoN8Za6IIK2
altY6rZJp7+jj0vde8HBonXU5Yj9DAtlEuv6+WnMT78284NhYwabi5PkZlyCd704r1uBh8ZdbHhA
0jsxn7qucujebwEvv6upLgaHfOVObOjTGAmUhLIqgegLAa+/j+7ER+5H+mY5CXZMze5HErt9Une7
KvKrdtkhHecHvMH8JOavK5IEVKsRnQtlLC8kWIawF2FjtNZtEDi7sNLL1D9Vhm7UcwclLNarzn3g
moI7CyMe6FOBK0+qGi9A0qZPRa00BtgAHi8Gyxpbrh0duksNdds4o4iEy1awu+D1BLm+TDKc6XBJ
CqINBFLMzxPw6j95fq5qCAs/nyEKquUeoHMAL0CJk4R9xsmwGufqSSDKzNnLWqzrIUZrg69CkHd0
sgXloPk2/oM1Uv6o+1quODtCrldcb/6FWqWB7rpmz1t8bUAvJ/oP2p7HuDkjV5Wiit7u1hl+qvME
qMTCBfGgEfp+EPCc5W4OR3N0gV1MgeuwmNWNODOrDPSrZ5diUPpKDhLOdQMQuKzPNzXXU0z1ifip
zybTv25OYVTbOpHKkXWKiqORYaxNHBVgU9ckpYpYXnxG6CjpA5/Ws+QgiTLzYliKS43wOwId/0xQ
dLixjTelbKLsx0rYFqoPTqW25HwKwNV5MgzsJJNknqWNPRqNXrDQNHXzhkTp9U+8INA4vprCkBRT
u5p47YiHKZaKUQwooXecqgyMb+L+RrohvLEm8l35bTi699UKkHZgiChqAhEXbQYvQjCG5jlTHBjT
aw5lbPYOq0SCDNbUV+0kQDDqT9V0JxMmzMi4iuGZdqtE2m58AsTKKKij0qUvq9vzjV8fI8ustlvh
+RF+3r3/kLUVPOpfSgQ5Lcacr6HptJsaNDyx1NiMNPEyVmWIWp1CKeF5GuxuTvXb/XHgpnjcJ04V
1ZzhR5xZ6pIe1cXdKw1sory6uWkwMES9IdPQf6g/M2lDRV9K9xbrlIFmbtGGS2B2ffWqjkNMVR9h
0ShgxSnPo2DnoFG1K0zMommzhK4NWs8d5SNID7xuVGQ064ovxWqShgiZu1ud2uYA8MF2LCtExZWC
gaTurTMg0ePxiVmCxaZ5KpgmWiJzMe/fi4FFE4ZCSUJoMDTRrX4eOdbwsWzKGzkm8AUVDZlm+dhD
yx3vvRSI0rMGHiXuE6sn7bhhTR83qinpw2EE3HZUe/9FuMuuke+9da/KAvn61othSDbzEt89T0VZ
D/iLBflviZwEwg3tOZDRgMMW4t6lu8uIPHoKcW1DHuVBZtz6jRrYr+ovFvSOfz+19zHPW2GSrCpe
y0hyCW5wondM1TIZ1HeTcR1mHam2kEfAMGNhmKAYeK0GNs2aHXrkXzMbDLCFL91lv3yHAOQtUgFF
GDh7Utw6oKRMMhFZi+m4lr3xQuDU1hUYmc49MTHfjjFmMY604V44I4lUnea7vRqys9fycxN91xKI
oHzABH7Mqf1xc1v8aDvlpSZ3T+oqd1uscw6x7Cl9tgI1js2LxCCsZz8MeW8n33NHX2SWppeNiiTd
HOqhhs44I8grz01/AxeGyRRLL/8z2STRjib46q0RgL5cux3lp3qS6VYsuV4jbic7H/tmspNBunF6
UhiAR3ecHMbcqOvj4yKFC++9XuU1kbnhGPC43+VJIKBsCIY/zBtBYKmcUj99lWzu9VOVpoDWUzNf
wm7FLV3G1fSVwO3Q//3a2xOYZagxFv73nzzUllVGqQQ32JUGbvRyvo/ErlyunUXEf7lPYYnETltz
cN7s+qQglCv6vvpJYqLPw2bKXiFiO9s7OAVXATJWC3hnMb/OPNz4qUmCZEO3hdw7tsHGcjQWiilY
bZlJKUJmzK7vmBRK4V1BkogRxApxyyypnCRdyrNowoEM9RyPq07FVfJMXvV6cEO3T+QSetFq+Ryu
5wp4b5vXP96Sej6BRZAPfuxIZWQmosqLUHgSMZyTwR6IJUo9SWMCBAcSPK2XiKWf+8lk5IAlEej1
UsgSZ/Ow9Q9Gt1MFfdDpGWzH4bojXPJpeC54OhXQ9ExTs97PleeZ7y1CqAxFlLzYxGPiByc4lJyA
VszCo+W8WNGxLVuWF2kViBRbjDmaX0qkjfSQ+uu1dkSQvbQnYkx9KhchTOodTeX4rs4d/KLlw1u5
hNzEaJS/HfbuOvcMKLpDRFVt+tQXoI+pxuhqWq/y8Xd1LXSh0C5IGAym+8mq20z1usYY9Sp8gYYF
SwbYH1cixBmmpRNAneYsbR6rfZgbjQ84Os/pnWY2qQl8CBjI+2qsRHHg9Yp+SmuBhRWHl+8Ohbbt
p9FdBpDefhX0Qut4i4ldGbQXludiCTZycbNtllyK7HBpDgBBqPH8PFXWHtL0PMTRpCZvMGo+t2jg
uDyVk1uhMIxYczm0gxw9yOzH/KMmKLvJQ0hu4zXegTfMEg6hzVDp/Ll6gkOk8coY/+b0NjL8jQx4
q88zkLwK1L9FQsr1idHLJmR8zII/lYYyMGQ4k5qMVrFReJRJozgtH2KQtbxqcFZXtxZ+yxeGPXJM
zq4/Lja7gK5ETI9zbVIht9yJM9di43H0myR1NDwDvYg+W69JkS7B+bbcuUIVa6dKidEM1HcZvAnS
KNcSI2gBegKNrEG4RLgRgzeUjBM4f1gOEpne45Ose9I7Wo302zov/4AbRj+2RZaKfuJTZWItADUW
euC37TtXdmewPMMAIaLtyf5CkUns7XI/BVqjz6oowEzIzm1/g5gn5CBLvS6zgUikMfrMRDVIMewr
ykksbyNs9CRd0bJPgLPDlO6SOzBIWyazOsnnxrZvrcXiVhV5T65Y3iIx659J+9Z0wRnAW6HDzuPy
+7xNljtFzhqLZPsTbcjJbxzRfUT9Iuy/rfGpzI7yO5CoGO95LlWZETX3IlDfr9ZjRUu77ooUuZny
MKVSNtWTuk4es9hGbzH59IunxfPO39iTFNDV+5EcrN0nEKTgdtH/4ZLfXqjxolGb6o8CUO97umB7
p5qSW8ERp8rx2WM7MV1aodkYlurSlAdV+jc6e2uPjb1eSZuSOxNiHec0THRl4Upo52Fw8o+WmKhO
kmX1WUccPT13pW/6uNYmKOhxWFztUqpRLDmYvG9UmL/HsoZf0BygTi1MMCNPptF2G+ng4jniU+oV
4WZ7Lzf0K8Ycaqvpy6a8t8yqCQTaQDi6kkhmwCh3rZYK6ApU3HwkBHgfyn7G6SaawnaabgEpEn44
EZ6oJV4l9vYqQAn7Fe3pWIj/USESIo5KVE+OFWX1e2oZmCg+qhNq8Gcqjpuyn/QtKMGytiSYiY8m
2+V7C/KOqnG0AsECU43s7a3e7HwuBdkXVZ4T4OI08o9p7HyZn04XEaJvOMipfVQWKQKRshfUAK0V
WwzW5osti2NmzrL3q8ArpgtIrN3Nsr0V9ZvEHmSYH8cxCEuMNzE0CR2f5MqP6lET9AHknVqmgBf8
UZdGwWKzxSV4qkT2WoUJ9ZcmakRb6Q7Ozr3tRoHIlMtVlcY1Rf95TtJXptfHcwKRayqGKhSHLeYU
HWSEnEzArQFoVmhOh6wyjc94XPabMI/OFlrfUd+faFFiY7lDeKqRPWlAdyFPT51ESh+3vIU9lgwv
pOlDmz6obwWNtvWna/ZRJHEsqrl7kV6JIaSSPSTihljd8jrkf/QkcKAu18f9aK9MAUKoOAt+n0hG
EuDiZe9YaGg87P9MpXQ6a/h7wYChgexSmAFBSrY7Op8xH/lzaLS3DGm82KsC1YQ6YPKG0BLjykNU
aANfOS1k2GEdRLlZn1Uj4bF6/dL0wZhGNzcFjARqmdetDCHgiD8i4cVrJC6EWEpIFq2Hj9UpRtph
0AzoAiyuyf4r1U6adQhUoiqZ5NUL8giQc7RUVJTTbUMK5aHy44ikjD/IVMvQPEyI2Qthelaq+KtU
9rGm43j8/3C2PjwhRDLHP3+9gNaOtiUFImYUFg+aptEQt7gbfwPZdfDADxBkXvnTH4NMGPk4yEc0
OAkJMq4yCMyDYRJgUmE0QEJDrk8sppFHZMs07u6qGrwXJ2aJRfTymWNDHiBgLZbjIFGO+JrZGwo9
aoFSZAX4cB0GU4xgCBZmm6zuqvj8jFzc0PBdHFshIBir8bR+s0xwzPn9a5GtxNV0GylyKkxr/uOe
JXWsHv7HuRlbbs3CoC7VwT0ykAhpMpSbfq+XG+Oz9lqlPR+aL6cAuJQCR6jVR3ZueMhBZHJ4k8ul
8ONS4O9uF8thMgXj9wmQZ2BI0kojfLXrdHEco7o3aYTxyv7bHe9fG5BHMGMKHnijKZnlK77EtOK7
s/ByRWfbVwhb7G55qXbJSzAhVrdLjIQYJlqCgp49I7mr5Wx0HIhBgQLksi6ajGBNSn9PB4pIKI6U
KW/u0Uv6OHAw5z+66+3Q8VcRhrGOImQqGz/VBd4Jzch3MFxTciZsZv7FTBFVkvhKZhRzeBAFtYpw
q1fP51uI5GYrmbsTMrXhIpvciv2NNIvqJh2beg97EpJ82y2M+IyslRp2aVq+jfuVhG95Xodeh++N
75zuj4vuvuD4ilDXUgNaLCWYwIWecM74X/eQK6j6LhTw1wM8L96mR0Eq+dPf548u5BPCnuXlYCRl
j888BCivfdf5ZWw+7YZJocIfbG9QV4Wyq+YnsuL4HCiT5olhe/5xEAp4ki619UqWA9haG58baN0/
zxogM888BfuF2MFOTzAFnqWlE/scUeE8460vZ6StGKY1WunPrVvOUXlQyb1i9Kx8McpeZGl9aqfF
sedq9lvtIQISKly3NijtpfReANqMKxZ6Wgim7U1Ii/J3gc9esYx/Z9vcfMvf4a0A3kTdQruDMzZb
Go6WdPzGKgzl0fOG5S9s/bIJrN58pkTsqdV/6b8OBSvDHHkFA+aoJxm9SUxdYE/ehkY6+vIv0opN
lFrnMoqMosdhUXK+0NepvhgfYUDeKleqOVR9StF0ZzcNU3vBjI2PsFTTdH1IdDpcLD/b8/wKxPlC
ohBRqyYuUB7DPSLVfu1K8qe1X/nI5AOVTLu0+M6QM9NAkhfQD2W4lTqH3wILfzM7AyRD2fmFISJZ
FGVUpyPSa4D6M5AkQnu/Y0ffXvpMxkb78JeVdhyzn+gEEYKVTxloqu2K/m8JWlRnWWr56x9KQjlp
P+V7pVBGv7njKb+l+xcJ8/kd7b1WH+PhnpVtbK1f3Aix/LqCVzX+3kvTtlhJUekDlT4E4cE0HzJS
J2ps+lBBDugJwnvV1U/IcvbJ6tAHZGwz1hzsDTsfZkp8ZkjMoWeC/qe01D7JFwwvP+bHTV7ScB4R
oOPnHMezYnvFsEg0VICqvt+wgAJtRmRkzW/xdkQhfg3UEJ9HYXcgjz6+K/ewQVJfjpiE90Ehzc7E
mjggn9gdsVrC31ti71ecahmd2tRgJYP3caAZKHAOKLM1nV0gxYBh022u3A8iVrEZOwHQrF9cOt4L
nc30QaShi5IvZVhbEO5KH2aK8QPyew1VlBYVy5WWC9IoSt/jzhnVkeJWP13o1bxgyMzlMYomV1k8
d3EwmVd9YOqO2X/n28sCVdwi9JSBvoUSTBftn2QmmhSqnCUBULKrjHMOnv9PZgcCjjBN/kYuKuf1
SftF+JXaBlxb/Co2d7eud++1Bf3eTuegx8RSq79cH6ktci0Qx0PyaUqnE20fGt4sn7XT5m8Xk8A5
mpM4/dRGUtTfeyyEv5yasRLrTaXfJioyc4R7vb/ekbCaL0qsvSgbtiVBD/vtvM4v/vwxRKXAY4lj
6pXKuJ+jd09QRGYeRr/nazTNj32BCfIN3aNu6j0JeH36H9PqWPFJgkdFRmhoROFRmxHPoG1IE7GR
m+wntpEGWEUIx7R8FK4hFjxv/pUsZRF1SO6JgMp0E96RkSBEXC5mVFsNIDmo1FPnYZ7KNwwMDw0N
cyqJ3f8ZBpzHSSNHq+jFGWBcrK2nXbLahzNvOGBpYdZyEQkasBvFQqZuCMLM2PvbUlco+P+GJsEF
+VmUk3AaIxSi8EtrTdaXhNfJJoJJVvTA+2Dt8XuRKi5P+bkDyRbNSYASLgWreC4qzhwSmeGAuu64
3ZWZbI7pbyb1Q8YZbgeeaukBo2V4V4CqzNatHQjkDHjKYc/UZzfLUaGk3VYDFJUnvo6aN1UwVhy+
ZSE/Z6vuFhBhZVxl0mbPFIxX8SOljf0m7RGQT4pIlgZh1U69ZDHGK3vhJ/nH720uQi5Zsjsf9puw
cGCijnWFeYr2OTeDDBBqWLQ5EOi5OTCGJfKASUKtWnxVKzAPBf6aIL6Ejo1IAgMQ7NUyR//hkMQH
Bwbadp4Dpj6lQsEZ1WGtyrWH6suepDY87VnAVOjYDnftnEB8B4oe5gGYsy0v8QpFLdfLsInZNrrq
/e2OtDhbE2IUF7/x07KFRAjwwJF1vDQeMKGXuiuonI/XxBcMO0WkrsssSfFFbogIrfPtD5AuOwP0
5RmdFDYR75LX7CrTTfkOecDzU8zkOsX3eXddq7zJJCfV9ofmTjysbcSloqzqBnLO8Pfqu8/Es3QX
JHK3uLilN8pxRwj0MxILRNzVay6UpebYxmVeZgZeZJGa+Yf460ZWkBwXJsOMgZUwmLU6Ee3PkEo+
uVyS+xmZ6bg8ao83yS8Pjq1jveYFEro6otT2P4SNJK9OzPW2/Yb9RrOxfAI+4PMd9DLo58KUHVny
e3W6N2EOkVu8UEeqaLpPqSoZBsOFxPeyal6JssZ+R6cYRZPobJE1Pm2xs3UuHRnRKA2SbBWJ09uT
VEGD6J5elqJl5EzbS7Syn8tBnVHSofPyWSP3N1sU8Z2LFYK3UT3WM311/dO2FYsVASPqQga/ttCd
mUkA0kQNWUJjbVpztAlspOGhkQPgS2FOU6i79HFXtu8z8PJAOob0Z1nwuDlZV8mqqAQwYVwkhJaD
Ngubx0SvFXYKoyEHp3ENfhlmsBIaksTN+NNyQ56jbmDjccZJbVN4CJzkUQeOlIxTI1t30Ux3xBb8
pE3Jx4LcsNXSkH0DyPWu3AWyOuMZTHEo86At9kenb8RfuvBpiA9hMcxZMrUPR37xa0KzHDK3dl6+
qtQo5e/YhYKPInY8DY1E3EoWO5fsrREDzOV/xru2tPZa6llcZgRtseh95DZmOUY8FYVF5UnNETK/
IV6c/WOW9bWn0vZ2VVwsYqSaldxz6k0iI3FZeEyIHEOBtvtGxepOLR9xxHIBuWDdQbLIosqXbOzq
3EEVkV/tII3M8zEmFuxgib1gswTR+ehz25e8sBjJi20mjBbeScSMet+rX2HRfT0r1gzXDG1SRRGP
wZ5C33DA7sNyIc5jC/WpsIxHIJIhyX1YFtFpuj7RWehQbqoUPN+HqOtn+na+YVT4sInPe3+Z7ujj
HJQtZiNekZV6zi9pYpqvp8o2WMjhpL3pIlcayB+okqVfXvepgficX2jxL1Ej4XYV+bi/+M/2z/60
1Ne8FeUypOyh4D3Yp/Reh0ykJ00YpvX7H6ur51cxoTOmzZEpvugUcxERGSJn72BJycAS9bsB4jC9
12dFU/EsCf54STYYA0omH//37yGSEyDronlv2PiMYU+BbB3PoCtATvoBJzFPa0QxzBjM0vTfFYya
CAFZ99ZFWMIruVJiLM1FTAa0wqWUHEKV44sJLH3D7kv1OVDu/whCx+V0e1jOR82hSmLUQpNScTFG
YKWz3DPy8CyASCExhcZVv0o/opsmIp12h8OoXPMWqO0mTimhcfO/rqDmKwrYtKc/XC3ODjJNjKzP
UuR05hzds4Wlo6XxmUEXQnI017y5Wj5vWbBzwX6wyEpJaNAYRTdKqiYGNisHPmENaN8oioAYNXKA
Vmcbzgd3W9GiCW5E2cy5zIV/4fVfZnMWyYQ5/xJ73gpjg56Z2L8y8+R5hR3vy6jZ4QM1LPKSQmIH
zQBRsQ4vJF1aJS/T717z/9f1wvYWHFCfKmYHF9AjMvZ7HsbXk9PGr6pXf0xWX2bBcDRrJZ2YtHnv
L8RFq8Ld5qhb+Twihs05A136XMygeRvDankenB1TGO1Zt7OLB14Fd3e5dk14Ooi36TeMG1rNTC/s
yswyjl9tGoJJFD6nUE1RR2E/hULgVoSKgE/YvO8PWtz49tEs6Qt+pDr96+LvOFKGQ9LSRNz9wrHe
f98Yc1Lx3D9TX7wunDU56FHAse0lHP1W+TB8jLtgRuhBP5khQGQmsx4JX240i6oH4GkJQp35r29u
h6kOYL+mgHY/ygCwCkKD5KX2ZF/4GsJD1aDa8Zf6nErXwPnyjgWgYV/gZPBgHwLkOIBdpw6+B/p0
w05g2eZVX5wua2j4WA4MYW+rqrxZorx3MuvrHbSBWiHeuonvjleCxRvAYHKJoivtg8emaj1GLuOp
7evcX8ycSBbECRsQkC+gY76MjW9xq44oBr8K05IjSTobA0UEuGGFaMPNCSq7xDPuJshEb4MchU84
CZeWIEVX5oBVqdlXHpT6mgzT3vxADyIg3XFm2HI0Ou5fYEbT7pAnlZ3YhvGFvbt1k3kpFFFTtmFR
MJwmDGCjLn5OaeUU/e+qqYjG9VOlg0bfbG0oNKBrcLaJ14z4Ntq97UMN/LUsR2uX8ejYrWybcl2U
7AGFkoJPFhvIaL/JJc1G5qDyea1FukMY/2T6cefcF4ATUrlTGdiPOXuUElgY1b3Ff+yrfGbbnpjh
piYRxLUE0uBw9/WBruOFaGzA7ygOktkHddTXR9Ul5lvyBLwrUJ58IS+jO1pBfavUlqg3ICgNVvc0
Qke19vjgKa9Et8/5ZTb0CzfVh9MosecaxY0IyYLota3BjTAk9//HJ4QsDjhs3QZeOTW7+usGHR3T
yURgVdKqUjXwuDc5EldoNaFqZ/b6JlzeZT7bgrNKJD+cnMG9Hilm7+Ry8fKFVKe8nWZ+cijwtx9/
XfLVVHiPlOJknLssWGzofI84KjbGp9el6ryVQXz8H9aOTER8lVPO7nNmL/eWg8ImYmBl5jCmNMfv
iBe69O3lI+CFyzCVa6SBellktY0cli7DB3Iu7CBQeYDFtAYYTPQKL5WCFBvP+UkJCRO9b1gqOXBX
jBgTz988kvCTPhV9ZmPwabz2OxOPifFZz0H+XKiMWhkKBnluoAIBKOIWg3NtMqn03wco6PzLyUGa
wH64wqLNxRTa8CA0mPww6UzcLEabC1eShloiQaiu5eTKCjpV3jm5dgDxIXddyvgsAzi0Z3YxpnRO
2qx3A6+bupcoOQO6xJlSe/kRphRSv9x0ysoftj6joRjMrILwppqRd8YyYpvwribQWS3Y9NMjPtth
vj8bQBOgRgjlFcvU5JSJqsvXZMqoN1UCRHcOFNRnHcNYVwWf0EqpRKoncl66Ri18C+xXDWdKOM/C
ZrtpW9WqJmieCdASloNSZIprwDaJ/xMQqDtIGf7rUBSXTMAGJwsfzcgsz/EzOayq2geXdgryPUWB
orpcWRCFWUdcYLtxciS4UGESCCMULSIu7/yWYPUT8VmF+zIgwKryq6Xr9wvpl87sWjN5T2vP3lrW
oDZF3Y+deba2W7rxoRmwtMa8SjypDKVaV01thn2BhUWAw/8g6FotirK2er4trnPAGJ9QeH4+iyWX
B9g9p4wvtibLrtThyjAUWtkVO9T0qZW9I/FgGf2Na8wjIp97dZDFUBk7mKc6DoO6MSmiwAINGzvV
d0quHSNRYqws61jmfNyBYstUDQrNIMFxr9nVLbTg0QztbVtmCyUgN26OQOCGp1+Q77zOw0Zizlq7
8beZ7CBo62JOQ7m/i7jjFQBMxhJXkbCa9m80s6/y0kvkY6p3Cjkcvs5cXlGiFDUS/B7HwDsoKKqc
6mjF7K3aNjaKG9btxQzkiD5w3fvWZlJnfkkLny23vbqWCC5pzgCYtgSR7SQyN7yAmIDYuq1ELpT6
i/T5zrSIN6puv7D+WMJfwRoSpNAIVHzX2WQHB22MNWitu530/LyDrKYUqzFXO0yLNvKSoBEzrh+L
MyekI9osFyqtBfqIcIBmxIPb2zB0KM/QyUNu8M4UQCvZdd3y8C8k6EKjtaN22NEzsfFbS4hqCtL0
EG73VLuwiPFK857FiRwVnVXpjgHY7I/hL9n4weV335AAbeYxcqHHhgEXKP+mUjdA4dchdMKlckRu
mxSBKS4gQvR+Wc8F5++GfaOFymRuLgdXxU7i1U9xydYlgVgQP24oaDr/ftj9kaR8izGuu5CSmVRf
pvvl11UjY0Rxa+xwNt1d5CBGYUrsgpjnDwHlXu6wWjQdxVLoQjOee72NLmRtcIViYU3ph5t3iFEp
C5P2AjBoDF4R9vLkRAX/tCdbKPxhNT19Wi3AVpy83nH9agfM4EUKLhJ1+x+sbyaCGZjd8vWJny+g
U4y3FKwPXF953++y9e1pPfPJsSMTd2XTZcatslAwKdGeDwMKwjKR0V8OiXgfzW1gJ6M92zRnWLVM
sWEKJ+NZIUf7KCuGxilFPn23TO0Vu2fEz9WEkv1rukYjJBRdxtSYtj42bMh+iMtuF9sIZ0JRWR3M
SbgoAxZ0JtetsukQ2jWhLRKMs5ydR8bd+giE58Pi4RqP32ARqBveiMB2NsjJJCJZnOivBJHNaZmQ
zzyo+Tk4hhEkE53AzU6Mqj8yyFMLsM3EVmW8DPp91oa2RqTGo9mlWRf1gxaCkBWPvwjrwVnydw7L
8Rk+v2ZDS6NhuzOBS4Y//Lbmnqevk+R3rSPlPUsLj3zmXGstbRgh3ryytCYfXPgLrIdBk+rn0TAi
bt6FPoonvD7kL8rddc/55EZmlRpjbe/Won/fJIW+fK3j0pzOIS7Fp8QvC/zTjTOMKxbSooUshmUv
pa7xLZZTT7vqauRGKs7A8W5DiouVCHoTFq0RLzgJfwG4ehhqv9N5UIUjLxN/YGq69H0vKWXCpKiP
NaRtTjejK+YfQ1DSjmBWMKQ5a5XD/WqAS0hjJTM9rUlPHwkiZrgCHG4yBG+FaoSGCdX+GGai719D
OKxsJ9j2L6It1Z94FEcR5lJFy/4QdoTTPb7gDj7+JCA5Th/7TuBLZzkds9TjZwRDE3iAJdOdLXw5
WvasDvh1sBnoX/9YP6kqKt4m59/LjIXYd3RdMPfmtAQobcaZKdZ1ZMGAUwoJef0C01zQUDXKF/ED
yvkQWmLglkesfl42voOmPuvmgNJZNRwMZ5ITW3bW/4qWPQG+hYzTXw1nqHC4tFjNJSV7a7WxefHY
k18cLs3xsJqyXPSgqr+k0U2jckrDnCTwf/uE9NAAkizX6zKOfW7i6j6C+LKDwz++IQF6eGoPN8z4
PX23rqk1E7yXiqCSnkgpyOWhQxe+Kg4ZiTMsH/KJTm9QLbqU9TqJvGcZeQ/RQiIpHCgW0oRsiv1r
jdrwUTkR2+E/TDFZXxPjsxnS8JyS9m3Jk/9aHGeKlW0bGKIeM2/WhWYheq2w0CL4mmEXBMcZfWxt
5agSWOrQEEoegHpZMQffoJjsBOAmMCVRsNLWx5M8q+1zuf2l/1PMs+E7QK95pT5xhgjSU6zd5hgp
KZw3/VuNil/XoJBHkErJEgfTNq+JyI6eH+cL7yT1ANzptFNnYqHmEQ4ff5B9dDGFoyxkFFv5KI+e
OtccaBVgviPqfQPlcli2jz4Xsge9JrxaHwFj1bE+ECQT4ENolA58evkLZfuWjLZBV26rI5BnYcY1
E+b742lwKrS13udiPxVaIlLUXw368xkqnAGzqHGBTvP/OnCdP6ew6HYxUbjz4oWpN9mcpmYz7Llf
7M8SbdgGhl9hDxJbZKkTtQ79OMkAP9DojkNmM8l+qHoqJITpYWWEJm8SySlzi6/LoYCHkhnzFgO8
X+L+9A1V2yHWhScrtrN9BIEWAryL8yFWfKfeXznqOtrbQXr8fR/8YIvr8qRfU2DgfZs+R6pkNNZa
nA/UMV8eknuaiUeW/OvgeTTdsDiJsKm5zOTA8EqOqmzul/LuNoYCCPZb32KuTLK2M6oPNqvQumKd
2mp9I589o/OdNhn1kXTkrF/NeOibzXie8kumsb+FmLo1pU+OtKtue32KC8AzIm646aQiPEZlNhw+
nRKpfThiwVv4mcxklY/Hp1FzZu5tCC1PAI85c7CT28UxcErQMgV2RxCgOlfEumVl6qqwhCWnrybk
aKQ0nwAg1Ga3og10sOjNNSgVyE3kE4a7xMhhNSK4XN7qb0nlYVGWP7qu3UFwgWJsud8QPO8Q5Z4y
uqa9AjvD0ZkOip98yClD3qm92kGDWYm9DqzM3cVtX20Ssfq1EY4isSp7bki1kkYmQ0gSRbpuIvHB
ChSk4Uvwo392TIezqeRE/FMdQC4iTvTsaR+t67mF6HoqpDU11MjEl3SqLjCR8d6gy1pr1UJqO1Lm
Ovi9wXDYrRnU126nn2UnkMCQqanW7NL9UgJExQWrPAN5GZZfwsltqojL34DSR/bS5DCmINjrAC8u
PyNh2ZbudTnUrQyVxn/Tswq7mRuf0VD3s7ro1r7VGmIPFDA4Yh8s2haUfo2ra/GvRD/hGCVDLitO
hgiv86wBDk1B7KfYohI3LwCM0qMXZJG9eckG25/OW+zdMUIvrwbKLd/5LZXDpo+d0OOmLv1tpMdH
8ZH7A04cjSme/ZJjTZ+D2y2txcoNq1gFx7x+E+fEyt3R8xLGxszZ1nBQWXmbOOqsaFut+cK4PbJC
kT5203HXD15UbE4Nnsqa4nU1dfzk/SNK5X4TkLLltbs0y2rlzKkZM2QLxGXIIhWOpUCEO+JKAXUX
B3hEL538al18c+J1T6A0SeMHvLdtvb3ip75wJy0yJR6BBVMbet7vJPz7+PJSvFLxgrcSVOyNuxEk
k7OZyoNcel4m+YeUV/AsIpiI7s134UgSTA47iljLpEMpsV1IP3/vG2P0/lp/u09QbNBJy6ZryVxL
apmEYQejoW3hLMKT8U7UH/9DmYaZc6ndvPbeeUEhrT5CcCJ+HkwkaFYDC/aA4AxhHU+FfeHdKBYL
PnwvB2YVpl6hQ0rYpYiEiIinSsEzc5dWlRU6etBVcSewrTLnUbXTp6JCItChur0rZtaAv5+z3Uov
a/2TI2z6k1yErsuWQUE2E6PCSymqHrlh4Z3GvVS8dPXUiGV1M5+xAOhCvpAZsu83ISbk1COJVY+5
nke0in09oWFIZTy4Ewt1+URcEsR2hgk/cQ2ca1UJu9bKWvHU64ttOpGsa57tNcS9nzQiw0hR8w1h
fefSiFgKf8+93YUVj/3DaueI//SI6+O0vrpDH7nSjEqrT5sdMGn8FoipbHoqSjudd62HOme4yIex
PtgA3fuaQk6U8IDPRrOeE7TvA7EuXcppVXMgU/tYaN6uJAayekkktob7DaM7iuAY59+tG6bmxEuy
lkFW//I9QyK7s61HLCFPigbrvnvBYL6qNpmlGCcKmTMLma8AukbEjxKV6RBhivzgU4KAwNz/JbgY
4zX2y8QHDe+87yTpD81uGsDFsdcVnNVrDkQqzTJwyaIU4BOulDaal+wMVDBqulY7PO/Tj85vwhUY
i7b5BsNGzWxD2o7O/9335MY4g6AFN6M5AloJbF8SAealztTwvNdz5aD3SKQkkjrnmPptK68iNB+n
oNNeD960lkHPlWZ5g1Whr0zmAh1IhZuKytYwZwjs8YuH+DvOHvWSNmN7I8Vxlo2MrXwlLkKRjlqy
+ZA3wAX7ogpF7poBrL3Ha1LnhUX0QXWrY+hESGRQzfzUYT6PLK16F319pWVH3t+4fIAsCix37AnU
18+/3UIVY2YNBDULS1pXDpkeEJq4iEGcg6kKdeDwUAKmMFdnjINW3qURY5SMsw1dU6Jcze59m38H
Gw1eItxNr6QWa1q4RXTZvSNLXGgNj1/EQseDgtlHLPRBXxm9yLNBFnwGxYk2OEwqwJQM/tKA3exp
Pf5jeoKWKEZIBQrUbJon2eCic5YJWoVRg4PqcaMO9YdlR8I3fjWVz7XUygfG+ceFnO3wzsyGzOyB
DXOHKWw2pKY49nxRgx4m84w1ot1LC4Q2kS2oYPfJTPlGKTH438iLTid8QlG3ALkhKk8aw4+s8waP
vq6DfzmERrQlzFCtnIwqtZS9Sx9M1LQ86moJY8P/ZBQBLWnlTZY6c6grU3ipIe0cdqdWd8O+S3gn
ycBHf0yMJbFUbqvIy0KmkDZkHMTkRMFM+pqU+zjFbbccYgnPvWyQXDb/nSPvlVcBu1cKKsF62Gs6
ipNPjo36M5L3/XJzrZGgsQnwiQhwFDm5ISf29oxe2KQRZdaWHm9ph5BYCbzXI0CD0wZOhVgEonGi
tR7zekDx0c/6giL0Sn+HL3R9FYf4iSRVlZZ8ijZB+Vu7HDhz8mYh+4mYMUncdW4cp3CZLJ/Wkv4o
yQVXkM+gF0SxzoLltAbTNyU/9LoxGnt7GUINEdmCAjC1iGe4RF/MAle5aOatH0A8vpPD+LZd7vLR
hM46aKRSBJPOY0NNHRTvhc0Q1RjjJHqkqoZ+jkA9KfuSiH92Prt6FpwAqygfeGL6Tt16PGBwYehy
4SGJ2Z8JT0/NF5dSBb5DWMQU0ru28R3lhqVWwGW/KEb3pPRfm2RtHYSOoIelI4TLTchag8XsK7Zu
qib8CgqVdBPEbzi/RUy2yTVKu1GRU8P620mcLC4Esg8hQA/BI2AJL2o+6eZhkJ+5SA/MNzFFAZdC
KkPcxlGDvAugsnwkszd2aaowcFAIsxqSePaQjcsiuruENg42oM9lXtLDBxlmQUFO9eSQ+CcZnR/h
3MAkY31Kvcdyb6sSRRvWs1wXKHZv6ggYQBC6VxVkhifTU+A7aCJda7YvwQ72wd7YAwZUlXHZTFqV
/sIfxmOw2RjEZHMPaRtzBwZAGN34AlQyfOym41VoPHZH89J4gbUXk4Z0JGzB84qLHsY0v1g6nD7D
kBQIugC7/g65OFgLqWgIe5uxh1aCwBF72Y7LPVFeQ5F1sRN8w7kSsNsQerpxgZ71U6wVX669+RA4
igD1p0l1UhrNkEts7wH+Hip/ty05T3fFaleHcDegNXXEX3BmZbv/JQEzbLi8M2mX5Fn8Ftp0tPj+
+5lnmXoaAcuj7rOeIddF5q9hCIWLiaqe8ThSkcjnd9mYugWOZo5BwJgCzFX441lXSpICGn0YqzAR
M0Uqr8KOxYc4qxteUYzlRnLHRcYgaOaYFVRltIXJq8qF1f2rKLgy/I6u9wU5TzqW7k3jW9OTdI5c
XtD1zzFWHO/6SFSoPNOKvt263zG6mldlEkq8O+wK02q0SYl5U+ZAwur9eT7SN8pGaukgMwwDTpBs
sEnAO8Q6qrc2TUC2nB45G9QBYrLdmtjUOprWycKCNmeCzH+BR9Bpd7WNUHeJBC39We9CGNmgDv0h
WDaWjOLvH9uqoXs6ACU8BWqu1a8NgiyELGZVwEPhCLpiMY5FHpcCMrVw7Xfcjs7fiv44/+6eSpck
rdxmWf+mPK6a2fwyzYmaFklFLfczDAM9lUwlkxB8SN8hx0CG+grdMVLLY2MpdPTsPCNk5AjCUd18
NFG1I3ZxpEEgYnWxmzi7mq8bqTGn59ry7ili60H2SWb65sPiWTE+a2j0TQ936vT45jTgw+OZJzFq
GXJT1m4JIYj3ZblHV3334JSQ9Y8CHFVM4XPKOWOTBt34Bab0h66zSawH7Xbzp3VZvVmmkiNmPwqU
knFGZTKBZUAZECuynebWPtr3kyNVWUCI9ZPoxIWsWj1OwVvby6lkTMP6gpRrrBg6QR5oJRxiWaYk
cEwc6iZlzl0ioNAQ2YLnB2QwhCBvEXz5PT4ova549hsUxDYsZXUUbqMitJkbdVPVbLWTz0PFAzOh
O1K1XyurhPLhsn8SN112zR5YD4oE+F/t2VuBp+SWn2+UCe6zegXiQN0+Iz6lukaavO7i+mGEM/kw
4s+KSPkmBIbkp5n0ZCM/te5AwdKdEHC9Uml2dnb3w11wSB2OwZ/4ZlLvBgHQwj5q+Hr6qUF9xemk
gAr9ixXk0kq+areT7LUW/ZJNOPnn1KQ4IHYf+PoF8b+7IUI1JanZvRWTJr0zI1rovzdtNhiYwtLK
xATmXY4eJ9/jU1+YAvis0GpoUk1TvYh3ZVrsoSVB7GXWdR+IuL5Q791YPk3SWL79dsEX9diQI/x7
U9HddVzXwfDkzD6lDDNSwNtL7lzkQ1WcYQ2/3w1eeujCG/Xih3bfweGkYhBoH1IeWaoC0QW78vCr
hauwX7X9eyPF41JDUhUiShZEBMeNbp338hAMjyhfWHT3PJyCEckJCiOsf6oOStDXL0WzUv9FmWIZ
i/AHag80+e0gaGRBk1fvIEp3ALQlZ2Fz1S5+yZAv5adiB0PNoKZ1LNxykS3bx+eiRcnwV7CY3nTb
VKtFgAyXOjm2d+eaPnpb4SZtGfuAgTnrSuFDXhAXNVyaJr4geeuDY/J878B1LWpvje3v1dtBWx/N
21MW9JZ+AUnxnP9FIYVSx+MpBmtB7pZ6q4xt6zRLjaddJcUXa4FB7cGlYKRQbW183fXgj3Hoaikz
hgD99vuy4W7wExyXWr/M+10XZyN3FI25TfU+5Kkh3JDEnE/JSU4ywYjm9Lb/BZ87BbbC5Gs7QJtt
HGvEAPW4obUVs8mI5Voi+OBrdBhLcd0pCeQobPU98ifIUwPCcJ0RZV0KsRjGw5qdKdG8FTCNSqOc
8+XOWje0zVtGyWZfOfgXAL5PPs6VP33uJOEDQ5JOOM9CJYoGMR/VWqefGMt74r8oHbcJKyHuD0Y/
sojLLjo+qwQcySCMaVVVY6dCbGnnd19SrTsZ8Y6mk7QNefFolALYwRd+JT9r8YhO9i7LD7ZqVUse
UdMrzkbdKuZI6r7jNlZf4h3twMREg5QjQ4oh/KR+2uAhUo72+NMfGbj4haatqwoDvHMswlokwyTV
Fhgx8LEj4hYN8cZOMnpRWiNzU3MST5IgH6sgwLRmQUq6Lhj1PqIsMOhivhUW7Oa+3ZGMMG/1r1ZF
dONQjWRpyesIv1swT6X7RKzsuTg5cgymVStmHJUXI6jSJUo1cspoG1xOWt3FaFI5C4uWhZT2IVV2
RPjFJoXy48ZfYxWrEABMH6YZPAezfpu60k/PA6V7QOMWIaGTVf6jba7HN3b7Omv15nSLbdcfGy1x
W3cIEC8azlHsq37FESUudBfIFrf8foig/9CPB9LgkIHoTrPwOMSdumZKTHz9LcQ/4bySDx5jt/eH
0e9Nx1B7YEzCgKF8BUBu2pInEekqINMWpTZDqw4OtjLXebpvsoYwJeTAlUbkGW2FoISnXM17LVfY
nU3eApTzEpMx3Ey4YxtBTtQViX5AwwR2SvVHBOFmW4BktGw5S5z+ZxeTgrmEhKoSyz/1QC/yTOR/
F4gKJ/UBxqUIuxebY6rM+jMGZdAAL+fkqSfrhFmm9hkJeK/IrcXcb+DZp5kAMwCPXGgDkemfJwwO
BHir3VNz4+sTvTbj6NloiIoZW5sLqbkwbzRntlHZ7A6IgqvQdJt1MzaRU8DVZDJT2t/6bUo27h4s
ITAsGMZ9AndkDOxVPQFkyfhXLj5LF8LrRs/JRhfoYQynZViMnrdPJfvvunrbZAtjqVcxKTUyPu6q
0nwA9dw8FUj9nsQ3mAMKBxeL0Ti3gQ3moSr7UzGQFTxFaik7Dx3GPEDXdgei4aR9GSPdLiGUjE07
OPy0mWeCt7+MwKvAMWgB5qwR75rCWz1HQg77Nkw33VNRgr/dHhCaTtpMoDQQPrFLembcDB7rfz0V
963Cq3TuBfJ0Uu2EMUTXbCej8IXHyl8iM8eafXL5C9rP5XSpmJnIV360UYiXQdsqk/c8gceY/6HD
90kKiTecV47ua29mDt7X9xDq5J6DMzA0Ofm+pTUXjEOua7yveXsc3Pkd/TvnlbrmN/jcTgGIT/Zs
wBMap34vsuvqNz+fev/IPdbAqlS/bFYtB8SatPS+66NGFUKQ5wpvfEOSZxL564u1qAq68sdM2ZaU
PCdxga3jPgHWWC/4+M3A4YQzE35HLl/XwXt1MN5iJCB/0SZhP3glZ39qPFITyfVfYTM6tSWtVNAd
4RqUXgKFsBVN1wTtWHrR7t6Lb+qCOhY/aJuud96Vocs3al1fHeVL1Iopa/zNRbCl93ZQcMstVG7t
8frAf1M39XchkqXEGI9uloINej1j4/FHQrziy8h5IjPd8ZuRkbfTfgNsFyDiWjR0GS9ZfI/rbBWA
saeGx3eldU3oEWdqSnK6cBdrTf62CblUmE4EE6WziZ2eN05fZr+Ky0zOEeusehCkG4ZzRpfzCeDe
E20Buoc8BP7cgOc5AAvddWzfkha+tSzWzn+Ay3IWfGCsJJHBu0NPys1jjQ2s56c5INj3rz6VW0oH
gGEcGcioiGDWEVdz6002HReobML7f1Dlmz+ObGpAAa/kJiYD5q3Jf+g2cL6aQJFpDguLilWX6+8K
PTsQdTYB/SEWmGiL/wIYn/TmNaVRtKQgZWDoaouaHPLJKmvxXF0yBvEKS8p6elc8ri/T1gZR+xEQ
/yQ5twu/r4OuGZ76t5LVwXisQyquu4hRHmZygN2/odCL+bMJ54/i4fiQHFGo4ddX6rSPqQmrqNJw
mqfjXrVhJEoEHwKalOmP5UOu2eBwfVFG6gw58HiBPEJTRN0ZLzudvN012RZBmc1GRmszCPcWpwwF
94frQsEulmDG2kOTqnsnLN8bdcAp4+LKf/4BVEtf48A9ZwwtgkrXJGUhAiPKbwDUHpcn9kkuYRVZ
PYmpjaNgGJm/kyTL8mY8ccLMTtywkG5Japnf2xP7zJ75NwZV3g+uXWnJWbMyQzp1/9WAxPoEgDQc
P1VlQy8ESQOGdc/h2Hjd+M1BsM+vJkBv6YrWh6AIqrU2fXDJYTBLnouqt8z/Gfphxi+70gp1hB9t
BMYO4BVlt8IGRBPlXdzT2dtvSmVq0/5TkusInIVqpIFDTgDm+WZ/vbhY/sKIZr5ImhXL74NDy2Iq
5hTT/cvOTc81NyGwNFu4hnOBbwk7q2qnGt2RnSW0dhN3mtx3Y+1IyKc5+aBapVBwS+dSc5JiOl6r
Xzg24jF7twgzv9keo9aiU4zsptjf0KD8P6hl60MB0t16BPWrXowBv9HzqVIHuGBl+ifFOwUOXV1I
7N2Ngo/cYrTGck4YEsQcv1bc2zPtkfKXFGJRUKWiqUevpbkuGcA4Jg9cxtWh1+mre78keLykH6ze
yeLcFOOQbdtDpuN9Bk7+KkkbRfRvAafph0wSZzO25uTuFqvqQbnMuARhmFDiU5wnV3NJBkKHIyM/
HW7lXUAlHxH3/FHoCmBSIbfPIsvgphADpWCntrx3uUQnQBn/CGQhFu9Sa+OSad0jqu8wV8kgjjCN
LilltYmhLDOEhJ/qNnBxwClTQQrK1Ayy6AjHMovjz1uht4+Xz4IUd5WDKMzCuejwD05mUa7RIbcV
XBZOFHuBDpKZgLWgtAeneVjTetBlm+yNRUT7RK1iYxXVodEUBtQQWgybKdksmyLuUVMfenygIRHW
hjnj9IqlvMz5AnhR5TF09tww4fpqUtDcSiy93pdTaS28HFYLORdO1vZKiDBe63vtQGPWKI9vkzTK
E+/Hs08iK1mUAzfzFnNJ0o7LHBJy8zCBKvGEI/fGY4I7MybWWf+hpuFlUZD9xRbbbBVU9xcK7yOJ
Kd/Pq1rMNkrRg3H2paL0nES2+rQa9ENOHNSy/E+/W11We7UOFq9UmVYKQTKHtgHd1KcGPd3YF5j3
RgFLjk3GocA++2CuQU3Bh1Ae4Ei3A33TdKoV7pdvnwpi1XCkcITTnfjS/6tDqc2aGOwqa7PLNVCD
/kpcRloH18XntJJ0X23D0kqyIvHn9x0zRStRm0TiNDaaUJQbms1kHOYfQGE050KwBda4+KrJlDvq
KwUdSvR32tjJAuvdoT1zcgR8AGfjqfFcGxlI1o4ASPKpYSBlpbLGNHlDZXpdbnE4KhodnL51denC
YpsMIny7BUZDaKvl47gWKbayjOg4Am4r7CN4RCXtlMVmC7cM3JzCS2HGSp/TMxFPV0JdX+/9yLX2
LHaIqF+4ZFTRg6y5heV3s0g0d08ByCpHzA/NJ8j6W1+8ODY78H2N/RDTOm0LpW+usBGgTDMvcpQD
5IxcuKNqmIw/6sWfc1SPfDaIg43jxLVERKXnkjmDQsF1nqxqnXTiDDSmZxIn5FZykizWaCV8Kft7
y+U+AJF0YKRLebinQ0mIHgJGnPj9bX+qJiINlKop9Nv5BZlHKVkQIAj9kctiSybERsLI00G4xDFG
JOrfx9eWpKPMgP/GeTU+LlflGJNVkKvrR+FMdPWo6xKf/UvQ6jxS9cmH441Ti0oveaZ5uRF0iQDy
0tSWcYVwnfFzepLSgyiHcklY4UNmNix/DGPRrEZ8wJA40w6o479x0G2+Y+sa7EO7H8bQ2SKEH6bt
F56Bafn96l70/A/YRUVvtwzdZKn0rDGl4WxglHtbKfHnq4967r+nf0m4RJXqvwn5dzUVIlg2DeHZ
+Iu7TVGbJflSuc/TWNIhkLOXB67QEEglBzFusMWV6/PZwIzTWQGGNeIhuaMK4dZUZImSlNa+y+MV
7dlDoWgnq7cap9zMvVrVdXHVuTqoXWdiLa0BPdf+A91eNUX7i30CDbCwxfpWPcBoDmZMJY7d9LM2
vsj/AUeMJZjnYZGYOZsglEVqZHQtO9F7HXlJLGPanYlz+Aiq4jAEC+GCc8kw1IlZDpf118FnTqMf
zH1Hmln0WlkU8ZWAH9kLA6o7rbGZmcjLlPyg6banokCrtWuKtvfHNJx94hgIpgYrLbFDifmzQa2K
eCHJ+z3m5aV0hY0c23xtPrQ32Y1LBnRmReXr4EOw/pfEKXPDWBhQcAtMym6ONY+E1o8bKDGnlmWU
Ps+pZhMPj/XCad+JfVnIUL9qXbY6nwgt2QplvJtEThOw9iflygCaOngGsUgANgb5Ot95EM2fGijU
tCk+ec65B6vrLYsO7iJiRuaF7Utp5GVcFXSrE7eTqOs5h7wdCov9RYJ7Mb+kkdW6nyIYHivet9S5
fkrPPz6WHYQIQSety9f1OlX5LHH+3JVxvVqii02hwft2en/VHHsV3ncZsWtgE84wLsbwTE00Nme3
NEzawY6H/9b6+xeU0AitwUa7eePIiXOWjh5bIfGMArXul6/it/lOdJKtPBOzTHvSYl74AvBEBpIt
NG3OqUWwCT16Zbuyvkjhj8MxfcLxVBR1kfUzjuNTWNRDsJElWVS0WTsMLxn9pLI9JK46WmmRqAsW
8Y47nlJluOl5CusO4R5XuYTHvAJX5pLzxAMT1JlHLRh7SeTeuAPqXCwzWnfdsmACG6NMl7Fj2NQV
8v4b3+wlb9Wkbx01AnOvoxmcBKROXNvNbKQMmP6btQDpx+bkbCM4+ZBbe8h18vtKqMjW/bn0AZoa
bbclgWHsCgKbv9IEwyvYRaiGz5RoxPODetfd3N2scEaUJ7vdd7mQDi0B0+6BzH0R7HqNsyjXFeij
S5L76fs+/ylzWQvKicL8fOEnHqab7/PdlIqFEuw621tR0UhdLm8S9u/TaS1sDMzoEMMziloW5ivE
cWEle690a3udHXnSdBwBInqN17wAhrpulDnBRtCEI5/NLptWd6aWpbQkWO4yxzadhQC8mFseIpaz
o2/RD0faAbt1UGNSGh1C2zTU/Tda3hAI+Z7PcizKVeSZGwk4vp0jI7VS757hAsnH0i3o21v94O3n
VftWIzVwGKuXNbzsyjXZ0HYIrMiJ8s9wS7tezTgrgMPB1OUbUFLDGC0z4qasgw8Buwcu0Z+4+3uv
sdMXQo5Gdnn80uJLfG8hBGvW378/cicEla6NAW1Iqei5rPJQJFJUA+vZQHCsmBVGjr9UDtleYX68
RoH8bDWycg6XVnWFl6jmvvWyadQLxPmDWETee+0Yat6voKIO3jNlcjO3ED1wLtYwKuEOeQCYTYhy
FVBrNJQejyggxYne2RMNGJuFKiYYYqfoe4eiUp4wI+bn8I3Td+Lv9joKuoCILcJWpbJN+gV+RZY/
mWhd7ma1SROPBqw12QAbfw6OFZMS5Bd5neyLoKLRA+MD2qCOuD3S3HXfd/u607AxSQYVctinKZUB
+gFz8kfMHbuJvj1HjF4jWEmLpFl+f0DMSgwNxEC24Ik++nVlsrQozuBk5Mb8tTvXx/puJ9x6AryT
+kj0XsYY42al+zppncDTCDQLdnPT2aP4e1FKFmpkOeWbzC0Y0EyxoPE7flb91wMEnoe6o582FxvQ
WCgKQxodKJqwhjTIN6kyYDy3jbWhHxz11fEfnRbgeoyX06b5GChVdmNPGggh6Q3SDj8aLCfQzcHh
r5Q1RAPqDZpv2JLHfH94TpUTwajwWtcPYtsXeMLBteSE3I7f6cB4GvsYmqH8uDjIgjrrLR0AWqaU
sODhgGHe4b3zIkdbzKpoR6OmPYMWHazysoCq/2ZomBwSVxG6hv1mUhnkYZgl4Nc4ABgQYmI9eI9F
lBPnJ/D32Fga3+pG2Zsezo9XD/11xnCtp9AmWimhZ6Q/SWxDZgz5wRWA1M66fgOPX0O1Us4dzXln
OM+TYy2OG7xZAWBnqB6FGxAvsHLDxse8AOUVPtpuvxWJsF00qGsFmGs8g5GibcXPaZy8iUU7+4ED
4NsoJCQrpAyNdWwuYfgmrZyRqyPOeJO7Kpe9JaTBo0JKY6Vt2tN7uVf0EyqKUaiM10WtGR4i9NiE
rkwtkpx5b95GowlMkBj7tk/0dTJG/rjk/Bn+BZiK0hDe/FLWBS3laGVzR4/aS34qmZyJAr9Ck1b6
TUaC4jXqYWIh6jJiMZzr7m3Fva0c6jRafvbcLM8xDhfNHa9zahgQSDiBB+Brd4z1dY7mKwZoPlo+
J4NgY45y1QYNHYWI7b5OzGEgK6Cr+DrzLIdof0KRncdFfkbSbd8c90U8EWeU0N8VYseW2oXZCEaj
aj7lchSsi3TGHaxjgn82Zb5VCBNDQAAIVIbIidKhy9JEdLvrLsEZNGOejizP+8R9AuCaUP0hf4Cr
2TxR/BauTNlvf7iA/iCdCfoOx35/1ngGLFErc+ZiE6Q/sKN9vzUfwgcsEwlmhazVykTouFgDQekT
DBbdjiN8sNPbAEETOzaoXR8LCaKS5iJ8lHVb4ZUM0SGDbZlI/pOUMrAMzYzVtJCfqtYOS37oBT00
9kfzyF4FUZZEi3uGfJslf1ReR/RHzEhLIfRV+1ppf5QUQsU6Vw7BSyv2SXSdO9YbP4O3M7IYoVQb
QDWm15wTxkUKsFe9fJf4UIqB12Vt3L3fPt7l2CZ0Hl2w8XKy+tt3VoehxcGq1YTMvy0cDoKOSG9G
cKdczsxRgbNEaCJesR7w3neAIhBf2hwVfBhPRBe5TqwWN/WlgbwqhCa/5WgyJTmVjwW0HU3Uvwby
t0Uw+vlJS+eKLZXKQgNhazKYVi8E+yHHVSpaI1nAczHl3t8TNTArI6BJZ3qeX1UScrHwaxXhhh80
5RgGf+pUooo4woWU7E2dfvNbLp/2j4Zyi6a526flIGrPZo2iHdgzb5OB1VCSqithq/jJdlEuka10
gWWtpjsDyqWfvUQQk71yRUeqfmw7X6MvHXTa7iX6SD8uv8ac2Au9NEb4tGjJ3fEDPqHvc9uoOPHT
M1p1nh+Jt/uJM0wuc2bbn4PV6q9amFzigq6jiehWiFDcrnFuDCBSIZOiDslN3IDFSEjSxDAQ5YU7
jS3ctASn1wAaRbcrbtDhA1X9VgHxi1hCm6SWVWudnckhEVreyoPbPNRglac0VvZ5KLpxm0vpakDW
fYaREb+j3ztDY0YRIUHqrotAxTekAFQ7STNhb/qHklQw6prt16cmgMFh1BmUpro2f8nm9B0MueaV
FK3ffX0OHfA8N1ukgkN/F6vn7Xm/SiCH0aWzk7596NF/cykf/eNger7+KhsCrC2R2w5TocZUZ29m
f3YtSBdDU6y2hjUXRDC2cpXykJmvwv5tU62RauewqMnObsgqF4pDTZ02e991UyLAhFSyJjwncl8M
mECcUdNgyAmvp9eiqoLXPY07jCG+Daa2WwrkURrJ1JorcFy87lCVcw49jIaFoKT2AtrI0OQnr6P+
Q6f7FGQNGGOTjtquRzzOQCCU2cVJyoaT1ljN1wLUCT/HlZCFeutfhghWfPOcwPFa3gGQcr0mxvGG
2yWI8KufGFYSW3VRypnd/wOAtl3CJyVZ/6evNay7Ec6vTjJXMM0cTjHqnjzfCGrf3Vm45v0zHUzd
pA4tW1507gOFyX5N62B9VTa626UXUyiC8omxJmfVZ5aARqavBZBXlDl+tCYVXUHhp+cafzM2DZ0I
EHG2T7JTE5nbR3noBcp6yQc/I5xc9YUOATGdfM9A8g+mValIhC6Stw6YimuDv+c/FCNKgAHGxuxT
ma7B8BfIdzsRv7C/UHeczJTkUJUJvtwUoCEvYaaLyvvI6QOknpzcCMw9Tnik8MvvUyheOCrV4VHF
iszWGVpEpz53nR5VicYn/8P5dLa0aetojQRZgoeyKoDd+UGiiEtk98YPaFD1M30ll4m6IHYKVRtg
FNBRDLTed7HKs9aGbkujoq3oNowAXCUHl0SjD2AaWQMvpj9RnBHDGTHcf+ls0FB3+T+Co+Hc2sWK
FIMEBoiHQGNihd8rPcw47ZfBjLywz3wy/aCy2JuXFnDy173tEVkl8+DiZ0AE+wm/xBEX9QGfngkb
pByspPclPmKuhse7k/XXulv9DxEAPYAzcCdPND9/u8bMdFCIr22+ZIP/s+x4WbBcp3SmVcUdWbe7
SUu6eOBzzuNqDRV7cugo7U8Vl+CqxlLcV3fw6+DLq4e5sXYxu8BCBCwE1a0ugvbE4vMR0g8L3QfV
uSp8eYylEgrZ8bUt/URHjnhgGvvudk6K3clE+ftGxHwuP5rKh5q7ZceET5q9Xj47+exIM8grn0qb
zANGNHno61SJ6p9iTseLJ6LRmvNvhgh1od2S1VIeFKfqMt7Ipkr1TlEzi+hGeb2AOIjBP2Kch3kc
iKhV9elah0KFEy5EoTgrL/qHwh8BLtrIHUzz/yQreFmxc99peQn4ccuS39S6oyADztU0vR1t3Sr6
CGVLFORy9tTVOQiFblFzkd6kZIJckEdrYeTxf9Qql1LKFEhqCJ70vFnLAEdSZfPCPbeYig9FFIWW
yGTu25Ba/X/PVLNtGZFi6zv2fr9R8rZQPkh+Ylf2kQYWUv+wr/JmmdulXPdsduvmqt8NvQKPjRfN
dUAJ2IX7t3jLtnS6yJ/AQvum6IIVOOPndKNiBDR2f2wDrylCoEOJcdmY+BO8eMGAFtLRrr/mqQpi
PQcbTVKsYqSOO5qlOPzSSDtuNOeXwCVyjP3rNfG2G+XLOhXXOn9qWE8oAGPmo5j4HNwf+GUAqoL1
CooeKoS5cwpazqb1t90zUFKjlTumUFRP6UO8kuYgyEum50d85+Sw8Qp+Xs5t3DjusdWSV5kpgiHc
MR0Ak5XhAfIGDBReffBZAwQdxfc05Hu3aC+caEoaSvg3nL5KZr02fWbvU/DG2n310O9gz1D+/wOm
GsA8Ui3XaY1Ml7oaF++wcpw3nq2avIKrsQGfoLCL0MlhR7Oll0fJdeS1CXFcboEWFQuAPsRfRkHt
rzE1tgQ2vknN5USIdnEHa0JNvwbTmh3olz+ZzHPIhuxCmd/cLHLa5H6ndn/Z98CqYw/uGWay8PGM
59/Qqoh469HL5xsh2xlfEPeyddHanmsptUrPPHEtUZpj/7ECJlexcCIRFzRxCQkN0FXpIU/djpEA
Q6iaRAN3cGNSGOffhJTurPXh+k53ieWV/9Dbp0y/eTIHnAU9zDTMnSc2ZesCRuAfRbgW3hxlKnpN
bKjm9RFh4KOtExHu6oJVrUTYSdZyPXdOyFH4Z/WLZxVe0gCeOJhZmj4ikUEu74gF4bPccCw/SuGI
jNP+DuPfbhorAjfpzJFIalPFJ/JKZe/GKOi0PCr56cOVCskbyUdu7kPoDsKiLsnri40t+PxqLDdB
iFo+f9zrNAsXXnF1D+7DycvHF92msH60ac0jBm2w4qLCn71BaUv8qeMGy2W8KHrE5zdbHQjvlytf
q9HFMO8iI5rsDW1iv2W3B5kYYiabUMEgVTsfU9eEnr8JakSGOpk2SeS10nYQq2CC08FowmpMICQj
UO7xg57ZuiJf7dBZHrP8OKmgJz3Ge4Qopofw6S5ezISxApaBK/6mj5+Uuu5N3MyisnOuFrABKSQh
BALFH/5bFH5J2kA6Y/wpnHGzoWZtXrzHajYL+cqjksfhGJEnMzOG+XpNVXSZJ3gTfcXAR140326m
8LnN13BmTTvIofqY6IPCG1g5Fh8EZbsM11YFHbn0+X0bJN1dI79EojZkEvZyMMBRXvFfi+KnY3W/
QlXPX6av8sSktH0Aek2zrVRH2BAiKmWOGYxM/nbgJGrzkqPYWbej6EYXGsbM3kh49dGD43yVXWUZ
neTagly1U59tbgPSJm1J3wib6EAPFCEtoj0ZgFM60xg+B8/dfQCpL5b2TFi5VzCWGMDXbW3REjkT
kopBF9yNeHg413kIGqcI68eJFTDkbnyWjtuuSjjYMAVT+YGRXAa3tSp5XdNrEl8UzsSZoXYIlIsH
F8f5SgvmIQAhrHky2GiKD4IDnzGbNPAufGQ7BGA8dEinGB0g3H+aMXq8xvcDBvohIfUAPpOE21uR
ZMND3bXLWXwMAMdnrq2PwdCXOurcGau8yC9OpY43jJpAKacv+E+RjadmGroda5bxgzvPJURHT6WH
FxrcIo8WwkGYQWWzGlLe3R4JoHPDuSUyLnJXx1m1AEriKWEqtqNzAqMSqmeRxfXYdBrNkCKsYlrI
wkoJmIi4fAX6f50tZTsiwDHHQd5+c0CJuks6vhTCuVdE6vbEa4wgqH+jH/4XJ660AXZZjL+KGlKK
f8yqoykS6KiU3bw3Ewhj7Sc4RYaqFRazMvPNuXWfr4AyAKVJmUqYsfIqGEQ7BpL7kt6HT4U0jpgc
ZiwmIX5lXootVSJhpO6R0Owpl2T99XgNR6bUXdaaeofkLAeFRu74VTm6X8+2oyR/y5u6Il4dDztm
1JfDEQ/3wnKqsCDZRIuL2OGajwgdO1ZtWKXVTrDMnICZ1RoTunHXEdUo2VrpXPeEP9CiZuqOeCWk
eflewgcPTUG5ukqR4o6j1PFd9mFMWcsZYmz4Se/IhUIM/HrwUCPMv05/yKYoTCZuWxlp2qJXYKVd
s7vz6jGS9/ibpi9vXenD7/9b7NLyoK3pRXe/X4TfeFFaBLU5BZF627YW4NWWX03ItlGY5yjqBCZY
YBv2KyK5X6sw3q1vqyTzlXY+OzEbx/jaHkA0MJHAzMhvQmVQUOPepHX0YRHSrzyUOVv81U/wLEc4
O18W1CGWWv7zwBmGqO0sG9/7SvVXnE7FH/04MAgHFkjI1PdmJiabnxS5yhKC5HaOFJecuN4+YzEj
UazopVscsSjUNUaAl9r0JjOreh4ibrakVOwgp1NsDhdUMbn0zptTwbHSBnwY3ZPRkSCGMQ1354VG
a5t2P2yvsJuqbI7fw0CMeg2d3d3HpkU4TJIgbrj3FsWYZ0O8m2CDD0lEnhAMyu+R1JuT30IwVW0x
3R4He46CD0Ghh/DCsOH5zEKLI2tJig6vgbVRh5fYnfvbPJlZe79QmG+w9XnDU5B3qjgwOeyZF7m8
J2OoDuWHJtwovxE4699Ih62HIhytQD5NRkH82JLdH9QhfBxLSZqQVERR7D9Ms0leDMTLlwxfgNFc
guXfhP5TT6747ZQwwIQdsxIIcJaP+zL/fwIIutUzojkTC40a9Q7JEBcSyzRuwI/4X+Uov10WVpIZ
tCvXwe8dWHmnGIfV6Oe3p7DfPd71yV034zrMnmcj8TGxfepqd0j3nyl/zfXkVEdynbt1KBFUBCQz
mElAMsFbN27sHz7kq+pNni9QexxFA+a+C/FIVP6l5Z9r5jOQt6CGEJHGBH1Ti1sqY8j9h7ZouZEl
lnCnIwqSfsZCvPrJiKbgfBw8pRHwTfn/mwQMWtfT9iAABDRlDdmWuKbUYRrtI1PjoXuCw4ttciK6
7++uPXo/lhYaQN3y47vI26eNqttdpS2oBr0FrLGatKrs0duam55+g5TFL1KIf1BVZVOXbr2P9moy
zakUfRsDInp1SCeAn6nxW1wymQpdLD8YatAXY0Q8CIXVUYRMRH9vYiUz+C+b9zm/9shMvfPuOuxj
wRct5YMqUbhbVogN4Kdsv136iUToWaclghsc01H5hqMsZoN/faBu2fnBaBXaAv1zb5BDQoIOV4tE
u9k34TkbHnPk6f1BRS/9lGZOOFZusVb6lDTWGCOY9nFpDPx7RlmZaZPxzFsP9tNEMviccGW5fu4S
BPHv8iFulUkJZWXQnsY/cio3vYhIYjL5/ZJy2Ss7Hmqp5mxvg6v6Yzuug9aYbzotTDJgpP7Imkzk
Xp0pyNSkvG6DNjlJoeZKNKABz4+iGTjonHwGH6wvDGa6i1O8lkFvdVD73/mdnNz/CCSH0LTw0bPP
PmTmWo5ygX5XB4H1jXIFEx5k2XZvz97F/49P3yZe0Dr7yNDzoQoewH5MisPive1yACmz2Xvs5u+r
Dvw92YKu6Jcgaln6VfEfTKp2IGrp36T8OXykKG3p5Ja2bIhFJhDWG/TjCdcBzZZt1K7iq1Umt3vB
d8SfRFzVPsTXCVrcwsyXp9cdf8e53+N3AKeliJHFq/nnXxD55D8a8aq+yj/s7aSqTzYwbnpaxH/M
OUbiFy6VlO0YBJTxEO4C73R/pdBV3s9Ld8dT2GrxrkeVu/vnU26UE4nPUUzySqmTQey2qc4iikLM
lz2FUEiKY+Hn6wF+5f7yGUAHjy3cuRAd9H2Vl63FS4g4ytN3Bfm8+B1bc3V3DzACAVX/A8+hcUwz
hsQfQgy0/zt05yc5oYaRen2nZcoGYZSWZ7o4GQcAY/NjSSj9xJlarSo53vGhujBzV+kycMavHwvr
hObsYnlUx/HNhmgThB2g+AmmLVy1Yonlu4MAVLJsxCEHYsFcM4AL9WnlMIrcmpGsi3HI57ZcNgsI
uE6q29cx+wSWjuvlG6SuFxPaSBpqM5WmW8H+uaNnqfG89kv+kFKONnIuDnFwlCjYHETRNklCDCT6
vs//PQ0ES1MqTRkwauHut3VoWfh95X2EV/GO0pwIbMKudm9IZ7zmQW7rcvxXENZK0rPBeMlaFgb0
cLpXh0pBvN8JiSIqZlTHVwdJiSU1ytHzITzfBFzS8pvu6X8s/gpxCl7XN9a6TUUqCJSKasMyWMko
QC4y1SS6bI5u6e0PFhW4rK9KdApbzP32ar9FKeZy4fWq78T1AOBluZKQ3ieMWtND/gCUOoLBaR94
kyDiYO85LgNkeJfGUDO8eeFewq21zJJRVW8jSQxWZLF51d0ESoaeJ5QKENtvNj7yi7UACQRmeNev
kTmdNuCg3cZF6dGooeInViwQkRPC669enbDegk14e2Fs0Pe/u/ldmJEvIxNGScLShQUGsgsEe8QC
a8ASFUZJzNEs3B8Y0Yh9ibGD9N+J8J4yHv/MpQEMOP+HjJbN9wOy4ANwegJx7vphqOHqNATM3FhW
U+QCCfvxbryrVWT9kkWrTsv4dEvFCgr9PPS04i+lUDoyXPEn19FDXrbSp+bkeUVYbkMmZjjFFC2x
X20xwAf6wEEXrRYHFz0aKZvQ2bFwS3PQ+K0im21xBh5vwGEYHRwuRP815jhMiNcuZR03yNk6SlEH
+ZGUzJZWNdQ3RIhrSJyJZ49Xyd5P+8MS4ooSNJb6wnMjL9Zj6jRvKz34zjRS4AhoZWJmK19+ari8
dtVm3NT9YosqiJ8hUcuHwrDZXVVHyut6YF+1lkYAQuJ5GwnGrv+k4YAbSVWLHbDJA411xT+3SC2R
sMf2LFCcFGRNCDI1m3CUvDIhaNQl8Bh+TrZmgoXyzoi3XhhhHlNDNWE1MEPkN1xCTxy2DXGvdCBy
EIXPFShKSoJI+6VeTe7WOCj68v7jpZA0vfb97WEFpUIm+4R2v04bMmSb+UlofeGji/sD55NF7xUY
JJ5Ddh4dKib43rNWnEtxAgZQ/3KA2HW42+0CDf56Zsk4ZNUBOdouKROWkGJ8FrJEzCWG0mmYud4f
UmuEfEi2H6uMjmH4CmZC2HGCn0DhLzJsjnoyxHHm1D92fg3KJlXpxJyfOeQpfsEbCpZbrmjFfCQt
bPHdckcZ5uTkWLRk4z37/dUOSpwp3r65ZzLNfPYkFIaVWoVyvOiIzs5t1oWFFeOsyPQtzARK3mAO
CzHqZzhNtfCVpm85in24+J1bEpE1L+Or+9A8xw+G0raczQfQe4zh51aCoeX5EM++ieKhZIY7Gu53
tAG0rVWKJsZfJyHD/zWifn8x+QrV5aKdFhAq6NUK0D65OcPmtGs7H2SZkt4h06ALXT8uccv6xxB8
Zw8kUMEc8k22PhcV/z6te751GHQihLlDeW5WVHhgDAlBG/xXbIYcSydWpU/VMkow5XDtmfrueqr2
IniahWvua4jV+z/MCEhEk4LXPDO3xf8JDbZ0ugNPFTJ/mHxZENv5/XVCaqE/LSo09GBxGPyn492h
ykJsBMecCWR4D0NtD7B7dEtaqoFLsvGm22/RbLtlLiiYbYpG3C0vgSmlCNOEr7LpRFGxo381/pVW
OK8h9PkgZCNlLY03q4Lz9QYRM5pW8UaMVYrWmYeAum4n+cmiUmmKu8amKLvJ9JDoImDb6J/OZX4S
AiRvNo8Vvzydu8gbIFm+/t0qkIENjGdb9vHxEP7HMAx8iV+/+cEHEQWEMKfc/y1WTnHOzcF4clk9
etHxVXXab4rACVUQaGh9kdx7luw1nK7iUiV7hIeuB5xSqfw1ALb9AVWweWiWRVlm7gKckomdE7Z6
F+0tvi3gTiZ5eEiyewiZmWqBFOplRcb3UY9ZlB6//SFDhtkdfzCeQ41zlbHPF3ahuz/QNxUXe9tb
NLCWL82GWkBnu3KGC8ke0/e2w0WrGCgXGoispZp9+yxpu8GnUEK+nIsozGPbeNN5mBRVqhof33mx
p8ei0N97/5xFslTE25shMTnuMr12b2yV0HrgM+FiddfFhpny2mvA8XV+/ncopJGifgWR6xL+KTn+
i9wBIjwweDk3+nx7OQg21J55LlB/VqRKZeaPhPvHGKUpBDevgPP0YWT4b0cT27FbZ51cl5U8Jp0g
alZg3+YKzRJzkBBfrdSl5V8D7BU8LIj0WZBPKc38iHEuGYpiD3TscMrDej6diCNdIUgKyXYP3Jbt
zBXyD2bUbwB7/kan0NQSv6p6asdPBsv60ZvSwYnv/2vzGKtnueeI1UnUAV1eRAO7LIq7KRxKDbYi
sezTdlYAj1Ad91sHrrnlcqYwCn/YDwh72Jg2G82KplAMHq8L0vz3hkmPrBItqd3G42jgtd3EACzS
Ml/VPad4pNE1zIoUjF3fvr2WNs5V6KHjpyIyrZnT5iT0EXMSiU99FsvGOYaRidShuldrTN/zIRY8
JYm6aEs7RQypkQDSY6DJBz68RA67x2i1X3tC2AkxNQKHTKwdHKnURU1a0eWO9OinGlf0rth9mG5H
gVAoi1DL0Z1IFGgmfl77khPWKVZ5YXjRxFlG2JdAkGw70CQMa7K8+fEuOFRHTuLBrDxrdqZAWSWU
joISTa4hLBZSL92lsed6c06qMuDxRhFMsWTBIFXeA48ptkIPiUwFCepB1rFppSjsafxYRTCFX6iB
NS0QeO4Kpu3mg/gXEZHL34ehSlBY4+Ja6BKmTsVeWvV8pdJYByVjvZU++ML9V8F3fYLfhrnD7GqN
+wsxnRSFJimscXvgCTgq1uY9UKaWTBgVQJ3qxpXN2mA+Gb79bp5T47Qep6aN2aTIo76pnql1qCU1
1IReGwBh9IYnAtpwjEjoFv2pBrVSl8THwL9rDAThwhHsiawFMGtKh1IapMHsN93YjVWHQEfEXD7V
q/oQxPWhuzQkFlGZc3Qd+Sod7cKasJrkxQafUvAAG6vTCZojdkE6O8Kuh3kcvPsS2MljpiL1DLU7
iUx5ll8/+1/1s4imIlo7cpxFmbpK3GWz3IzoEF7KB3L9CSOJlrAvgDa44ebzTxBrJ+/FbGUGNgSg
up1gUc3NxUPfUYBwRHqCaq+tfPvYqKcfSemMd2Xk0YMqsVZsd7wo3DHYchP7M2Fzi832+l2Lnp1a
vBjmMKgEZIHRDKwLSgmO0owoPDjOpLO458zbMpVacEf6R+NxYJ8kR5bBiV76wI3h51hRf/u6nNFP
/d4oihhICw43xzlJ4+qwIBvWb8amsVEwvrORHcnNaU+rXcbZCQnvNrBliQO4ALYTY4OKTcIkyXiN
fLl5OjTM2NxgoapeDNJ3dFywW/t0fjemIIyv8/hRfDyfAn1gdpp3UCeqfZXhbksCXiLpqub/2h/a
oQNLJ334wIIJj9v7CQnG94UmI5BEcIY9VW0VPdldvlfAxJpO5OXzSCYkVuIWPvmVZmKV1rbMacRf
ibCHZesnHEw2DTTmgIzsmHIh8ywCYNpYeVdYxiWMTuwjjjFK1djHKTulvlUSEsVjvgxvDd7iHcDM
PKT0yi+S72gW5gNCHaR42s7UPBP3LlHQS/R41QrSjnAr6lPHW6VrvTkPih/VqD4aIXuN8io1R6hD
tuVV/5nXq1fl6qKQQiSRO6a8GWUXw2Pawm8DvkGuUBMH+6nL18j3CnH3bqh36X40j1ib0/9WnJLe
l8SPtt8kaMPXC6A7fOfN3iy14TATDVfnT9Mgf/WJ9pP3YhHC4t9S6vCKfNcf/JRilmGZLcQne38t
zfCqh8VTchU/9UwfNE7/YbxN9nxavQ0tE6NHxT8fTJhznMCB2PcHpjTHPQPWNJJXDj5ssCASajmc
rPb5gs3As7shddv/6HeS3IOFftFKJYt4S7q86wsNtrwUqUrhwZt400SjeuVBXmTAnqqx1jMlezp8
YX/LWAG54xhQ+QNIwymxgoZY2SFgilixfYsIQ6yQ7t9qfxqZ2i3zxnXZ+IysOpIl5Fy94dESZ894
AD+LY9V4901Fvqw/GkIXMNUWq3Wad4n1IOyUPbTz+1yqXooxFRKj8qeRsj1KPNNcC+kJGAJxPYqg
24Q6pFiqrt4hsJR+NEHdhqquBhUT3yN6AB75wA1jiTZ8LH1yyxjv0YkZKYmv92t1j40izSFCtg6i
1E+Gnnc9ppIYtXfXkoYfMZIN5t29AIVfJbNQNDeoQ4NCe54Du6xc2djMlBCJy8lD0/25qWkPz2to
bw7tMkVQD5uMCvQdbocRfVDARqDIr/Y2UQcf+Iq5+EOJOn1OccDuEep4+laKSzUcPQSOEFMVKKkk
tovz8Ga7BmQ+yywZesYWpccYrzoZVWJzhmE+8ZZc54Mk8N8bjUS25Zb8W+CPciXBQ0K+ggcF1x9M
YnOtIZ7s72zI748hcoia+iHbaq+l2Dq5iBp/NJsSqOn4yWUmukl9C7FziytS2+7CEcyfxoYwInl1
8gbc663KtJfsmUY5cBuk9Cm1kqseCRxgujggGfgnEb2Pl3uBeQfTPqZjLo/h71tYbinyKeeH/rGk
Itp7raiGl22oExj/BeAP4WRBTu2+e3kBRSBRrqtq08fmLNMYimbFL54KCO9Ui0UMPRioKAtgpvGP
cWGTceeKrUyac2EiVAHYSyQeDHae8viPAfNNtSA8llqg6m1R8JzR5Ed62IKuo9gw4YrJmp4l3LL0
YH7M/3bjuCOcJ33inzINkmNRwzrV6nDxiG5qyMbxuj4m2kJDBsbvz+QyNYOnvCKVcKir491yLtUn
0U9XJu1XVqrjhoiVr7o1q+3MRgPj+5HDE/vsQRLo7PPZi59pN2k2CU0vLcNyN3hy9VNCWc8VH8a+
sL2vB/jgdfHw3tV4GJBKHhmtmiatxH+tO2l2bBmERDEPmxHFbhGWurCTxyUvv+agcWApg53JSw6e
jUWfBdqssAicjoemOU5ejt8WqeWwSqfzOJ2iX9eMDnTdjPuK6q8C4eT/vsZVbpRTbzsrSgk8ewmF
BzXms6jpezIPrpSdMAC4RSsQQ8pe2/VwxTV3hPgCi9KbffCODX0KbCpuZznHh8cayQgV6aSewMAR
WVg+ikDpaLwt0bYVnCipPW4mDCNpy+RdSGUvxtfow1rMf+vfLSbNBxD1gi8+qEWv/14eHeFKdsKk
FAZoIZEAskgpe73oYY2tiQUqlAzhT+I3EF9/ub+NMO/Ji2zb4z5vmG+qfDLSN1dmZwXvsV+ThGNy
dhyGBHlUKo/g2OB2002u8g+ghGt/LFIbN1AUY6OkxS2CoTlQA8WALf1UIccb/ji/CKojS7S65clb
dyBAwXlZx0IbP+9Mw8HeNITWpV3XFUpmfBMTGj5swznJEITuf3sWO6ybsM+/cIl1q0h82NDNAme/
MDhkP8o3Kb5od698O2Jyx08lvkiQ4EBBjfdrDauDLru+Dse8nDT5dkhzNfWdk8iZmLIpJYpb43PW
e22J2JVKoAWiSnO4thUEnZRH0Lr7LlLRjAes+R3mqKicbGJ4n2fHe6gzTCDDodjhdMEK7FqV2oAL
9tpPUKMNToT5/qcGfmMFElhUD4ov5jmQUrxO1/C/Bbj3SVfzOB0FZywyLg7+4M6F6KNjXNteEiGO
vQr3hQErANFKEiehOiuk5GD0Vg0oOFnG6oWOvjXYXW3azjVXD9IKDvNv51SpY9DwEUfwa3fdt4W7
QQRCpOmzkV8Lf2YQtnMahszIx+B5FJvVmiXo554THMQiXXfsV1ReMdIq9OIvNqzecJQYvdl2rYDw
GGOhS/vquizrJcFrrMphh8MFuXwzZYZfX2d/Tvqts0kLLBS/HFIpjkb6RfIuSoz8ll8W3iMLDVEn
uOa93pXx0+mr0kHOS5FUeyJBPKDf7mwJx0yJhYSECBja7I3vOOQzLhqMq5L0yG1HAme1GHmmfINi
SEkTl1fZyvze2BJsjVyI2dKoQnLvscUqxaV6vNPgVPKfdZeNdJDYAkwu7CmCS0c0CqLDcjTA9dQ1
OQNKyZm/YurtjV0HZFYyfiFU3ZeC9NKzOoKzX2dlF5mFNj9Iujj5CzJW7ET8ouKDNixQnGZOFTSw
WJJkY2ogB0ONnFUD7KOMv6xf1eDhKi4pxqs01qVR0XGYWUYIn3VeLZh9G1MBprJ9VpgDy3Gn4p+7
Os6IGUPoLcC2m6ra3FipqMDL39eyIQEokuI7RLnz7CKezdxaBBqFkyMy+vIRe9fJos5Hq3kjkIhq
5pVD/KLPtZAcowPoXH6v7OBMvjiSYtdMBn1BtPVoN/+XW7NR2DBAwfSjd/s/a81Tslaf4jcGFR2j
AYlJqyDIj49Ppp9OWCIQ3rz8WPLUliGKdu7hx5bYnpCLoBkcS97sW0cVChCPuRjOe2eYQSTuvZ7V
4cYa79qBq9umIaxC0mvx0AZwCUGr5J4FiLU0n3xhX760okSRcwsqGJebhJ0Ko2OFV3sYn/16qGk7
RMYmPs8P0OKPR5H4iXGhE9rg161fVPdEcdrXjvXFPov3LJCQ9OjU7B72u9/Wp+2njjpUO5ztuffc
qwcL687BxZDwv4AZ52jYoPWJTka3nBQrKRbodoSwU4mjNH1ns8Sm7Fgitpqcr1dKXplndg614RIz
V0CKAlQqglIvDA5b/huCLmrcnpF4iOV7CO6R9ZNtUbFc6rA17+P/vT7yav5DFznojIpIdHAMNHH3
gzBGozlp/yUc4HLAjCi4j2e8B8CoGaTMv+U48LaGlaTo9OhOiPZOeCaI/0+B/i4ntC+pGPZCJKph
VvRm4QfaN4ZgHa67GmTePGMJxE5XdXGh1A7apOGxbXsqQz+XE+kLCuGDNzKEjes0PXCXcaHDgUyG
bmHV0gkq5W6hanaPiybTC1kCztetSd9JLui9NlNuQaI8aN65QyKIFXRwXVKt+GOcX30lqKHoCV7c
0C7mjiKYJr0rZMfoU3NWF11sFdiK/rkr0n73vizier+gnfwh5Ib6bhzPoA2kCq8wLsjtcVeAKaKb
7I4mfdcCAdMgLlDfiUf9xBtBZwHLQbB+hJa5CZhO61p5mm1B98rDZKoW5MJlvXWiCZB02cie6XAh
TyyyC+s2g4G4CmhuYh5sgMmvbtwiOniEDbqSNOCwVYh5w5lIo2ufBWKXTPOilHDxOxOHp04DWv4z
ZUFNubmnJ44DdEtF5/G3OHnua5hpKQ3MNNxDDfr9DCewEzMYJUS1Mz/ejsERYUlBqnpAiH6ZjtSh
SBAw61vRJLqZlhN294kTDqXU8TlBkM7KzP3wfBlIS3EGuk3ZdaefjRUkQsJfVX2P/0/z58/HMj/s
2JxLdr9UNvqwCokh0DRi/156y21Y/U54kwDoCmnUvCB61+4KypBViJRTMGMYPkqfU5sfmE+sMBb5
XLGLWQYWmlY4kdQf/r77gTKyU1qLg3OPj2hM+BHAPantDUbxMLyc5m250b6A64NL+j/OWNuT5x1+
Kb2lcvxZVaBX3K3ZEda4s/DhZV6hr5pdMvUTRUXeMC3FC6lrFraOR95lWjwtdvzjqcS4i0QeBtSx
DKVAxaVt3+k3yuW1n9k+18OoAdkux0enn8Vn13rsmLkqYMXO/m2cq1zOI1yuYW3VhcxiLYBafH6A
IrQvYKkqRNJBvu6ZvTNJFbSukdhmlrVtU7mh3N9DiV7sc388aFpICSc7Qjs40kcgmIFE9ceAUrv1
VxiO124K0+mvBZRjAprJkJk8HMpqKePuEoHW7DHvTe2OR9LkOoNmdC6PiD3MFTf1VnxkVlW2qJ+n
DkggjC5x96OrTtBweGNWn51MO5sx8s+M7GNE1bXyBfBaxyaIg6Z+nZH/iSFyOYGkul1JXTpJtaJM
KZMzikQPN5uacGNdle/IB3Yb86uEUOMwhaSgJxQu/FT9+aNJSVLL6Slc0a6apCm8gJ7k2WwXB27W
CdO/YorriwSWbsyzxQ2ikDgkQcLrBgvKvj1wVt/8UKfq1T/tXqaz1z21BMHXp569oeStPi8RUhAH
f0IJtbEgO2NTSOFgC2a7A5+9d1cTjYcNMBC9eyrXb6ZmqlBeDEGGwD+S1qoahyKqY7cVgRaTkdbM
Hf9JdlHzubY/3cm7D6BUG/zl448MPC917fcSvcvmPY7aS+rzYdp+8m66X1SKpzuzlDr3vrQ6Emzg
/mDQZ87VgWidU1k15xYdP9CZyUFEIJ+btbnyPMUrQy0aqMLY5euuILU3wAixSfb7w8XmkEuGej6U
TLGfMz6TYLry+gp9RDCVF/g9uDe/JLAZgddGpPz7QzTIssNUmCHmWPaO5JSWizEy8tQ/pUU7F6Ik
ZRG1vgySF7UO4AzwK1pKzwSE42TTffGxvc6VxnGq+kE5aJzeL6LF3c8XhH/Hvv+ZGq0yzVMhk5fa
OgZcqWoIR/Y7z8J6aqjLj2kQzSyUuHffHgSt0URRPTtjZpaCs79u6NdiecyD+VsVAXvG4zOL4U5y
QxPT/vo9Y1sfawBvySfZai0/G5P2J2Zbq9ghVAn9j0qHy+zhUjnAQ5ka0S/VgWBWTGZjjyciCO8y
umYWHQdptR22i1iOKRww8zxSWDecE39hkI94OvPOgLNFtTBGdpD7sLpTXVckycCPcGsUbp66e3V7
8LBG3Fh8eg/O+TF2av7tfeBvezJp88NrppQuRn9jQpnMm14e6t9kzJugNmA23HLyBHCew8h4PuVl
zDQjpD+hCQRCSCrZRoyasUCdPHCzisLGpjwZtqSZ+XB8w2D29MqO6YmA/eVI/+IqHS+1sUyhMXXH
te4RnJto/Ii7CwuuKmKKw0B4wHBBIH7BpYIC0gtosiATUlqXK1jXu2ejGhD/0Th0LKUWbSAVcDqn
qftnNj2kvakRBP2fJ4utwjXXGsBiabATCrfjDxhhFrq80PqDJo9QCCovCVB4WbJChm57APLeOeTJ
dWJQmLCwpV7OBkuE6DsoUnxmO2JdJu64P8PpUJirtrhgU8FLOTNUu3+ESm3ql1EkEk/LKjgOV/L8
fHykvUzL885r0untuU9DaVdH6QESgzbG0Cc0AfHwWlZLxDQX9zXCBqS/m/7cRArc7VONEd2pf0Nz
ySnlJaYgtd5gyd3sQ+Z35Nh3oUVLJdIgxGIFBhwgJCiPPjXsSvLxXWChlxMTwc0ZSQkUpO4VXuZi
8sT2F/qkVL15W0MZTuB1ZrcaMNAFVkkeNwGhPwBmuCTpDVCDrKza35yOFXxGhuPFO9zRs6Z5Zp2G
2c2YIWV3AQnFXQGPnQQUCIF1JqJtkS8tjNEmf5Zu9m8Wa+pT7J/QgDfKnS0Yv0EBRnEB4AV0IIKJ
7IjbIK8iMpui1aZYf2CFUU8ouAk/uCR08kJLBtelQYeDGcuD6sYeTwUaFxYw9u2Of2zYVQcj1eGx
WQpzsSbpfsqH2UCYRp/Kv2NlvNV+/p1p9xK0R+XrRoES8zHk/He5uwEPJKbzYfUsTX8ZqvfMowSQ
4K6tFdkZcEEptdouVRFXUYQRHN/vQXYu+m/m+KpK+xlL040O7AGtyFoXav07qISQcMhzm2g0yg/N
BVSSWFCR+fM9GDdyVRjNhG0bSKfveMONE5wZe/q9KzSgl1fLiYEQkUcbj4rz+RGvpkH3C3cq6qkk
ayifNNVffczJO/gujxlP3zKOdHOZJ4mOkWtN5fwipQam3bMHQCUEufvhdlbL9ckjS9IBXNY/kIsg
UHqOVLNIayv4Y3eFbuLhur67tnl7MDGXioUjQ3jv6c1JEF3nUO/c9wQER7aDTQL57gu1PD18bicX
RSR8cJfc6AdbzY3c2Jonw2a4TnHL6vFunhDoqi4RPpL5OSgvA0qzz4ci8tktzpj9vmASbnyvFq7x
qBjX1WS4jROt1Pp6v3XkutWqP3GABvKYjYr09Y55XsPX7/QPsps3czpn4OBbWjE97351VHGfn0rW
tbAT8iqvnIHaG9p1jnChZoaSYkBBofaNyqVRSyeK1Usx4V7pYVTW2eujfYCAZVjWLW9F5w8SAPmy
ZAF6uUASRV4D5zPuY5mk72LmevcccOoldvvxmsL4N2oZoMjFwQEMhbOqpa1kBBKwrnzaWd4MFNEw
+z5FrFuSzKA8CHWpWN/b98TX+EPNkgn7ayBeJx3IPgSz1Hh86B5PoZNwCG3XIYt9UL/GvG98Tv1s
osQbgKJsW5Bw00TDOXSq2MTpLjcJNxhDpAaPu6o8k5UH3LhLP6G//ZmGnTlJ52IW3Lb17xwrpPrx
urCw0XPOQzE7x35gUauhEF5PRcF09zBwdYzeyrnw+aLsdbnAVnrlYxjG9Wk3dgFJT/s7YLbEUO6q
viazyxGxXgM8VS0kOt46goBXI/BWGMVJ0AJUAC4CT9aymq75vHffJyFRPYoehujRqsTh4dOmpfWe
+DnlumS46tRMSHlC5v6PrxqwnfZb895bDFNhiY5o0i8dM4kCdGJjsD0CtRAXyfgQmHPWCvGytR7E
fJ+/GCxu0heq5GSyI3NfntQ8noIuT08NMfZUKDkFLo7vO3oMdijCyvY47AcDpJ3GTC6+QYl6W6PF
IDvxWA1VAk9Zt2aByT/cYi8kyoiLZTyXtrMp/llI1sjpwwjLoEUV2dav2LsDcHuj/+sPuphWP2J6
E9ofeVZUYhFj+FKuMlP65uome5vNewlcc194EAnWOwOhY6RzmxY6TaKM74VsTH6KjIYumHRAUdnj
sDriifawnBIMV+CUoXRtGBWRFIE/BzsAdJygrmZF0sQAFIzTFaLqCIIAcZ1eOy1Ywarl8TQInCWd
IH48PX/mcvgsL5dkwiU9M/DUjvQ5ucfu+xKjOxqugE6e+rKpXnMjkfcrY8vi0EgNrAL6hbOtPxxk
D3WPtb5hvbIBiuEQ48rGxUzCM3OD0N4d+Ss2sCouYXNAmUu1KvE0upBDBHWWRkKnB6C5/IMAs1Rn
QHme0+XlAI4hdnfkn5UB1wGef8ydeCQ7LqWPNve1iQvdT+1uaLtjwMbaODMcMSQjm83Gd1Y+rRao
noqDd5BzbcbPnlMW6FON+dken72idGbjt4ZVzDTl7BEusN+a+1AMXdgZFHLlXTrm9rFIsn3ktu1X
G792F4wZJVV1AzfkcbAzqQBDBW8eP4kT9b63rNJ4JlnN5qsCH+BkBd7yJIY+skO7V5Qpp/UOfyvx
8FdHCE5B6oPaHjwGBsSn3ucXSgvnUkFa9qjm8m6Huyj3Fzrb6KMhorQ0ahfCQ9QdzC4uo7alAsEB
GTmz3vSeKoLZhcCidG5MBSXrBmhzTq4XrnZJ8rc8ZUeBA/puRMyNG8k2oYxc2R05rhNA3t5uryOH
PfRap0/HEmNUh21DH35kyN2fnHcYFWHXiAjzZVkh6MOrGGHPe7NB27HC5Wd87x0kTvo+x2pj7vjO
hQ1Hc1cK2zdyHfQyapuniR0sCSS5RKUgNCQT29igtKXL/vnPwwv7dpPRszNu2nJYxkOsuCJe4RfN
D5aWXj/OsOv1dJLN0hmEGxbOscqtWQipIA5M+uTpf1mllV9NhcW0lO3gs1eyc2IF2M23iyI1vdR5
b2P3yrkuTyBEWuHds/RycQ4QrNUdYvS5WgAvlKVGG3TXhjxnNtd5DiC59qpR0biI2MhnYUCd2Vb7
FLQRNu4y4kxI7Fcq1Mf+HAwIC2pLLD7aeq+yHfl+b7XsRHpaUKNk1zQFmfbm95j5OUTAtWQTOAqx
CB3hnLAMz/ltr0265EiULjsEjGPd64uYaT5dFIOWQEAOUX82TmWy04zp/4RJI/RGGXEXQaIEWk/9
N1bodiuoJ8y/HKeXh/oZ91o6hj0Otwaq2kgMgJSod0O1fXYIrd53H2MkTbKHOYSZqiJMkKEB3kZ5
WBZoTj4+ijmtc2rnTvwgbfO9wGzWJvkWHvqGlXsQDPe691+rkGz8jScX3YKZ+EGspC9iJCciIoAb
eRw1oCfVZ61kJNS7ja8V4TlsO608ms0Yqx20SVZu6Grhi4AZ1PrM9x9CfejiTiS3Awv4CqvAC6pX
+in/TNJOCKh1b65RVfb91eHGVeJsfPoUb4L9eSgYUQ7zIkTDdbVr+pukY5OedxTEuJmvQNs8CozL
fnLLAher9YbnmdFUKpirKbewFHaq+ZF3FVvZkI6pjPUl4tj6uoNh2/1fcG0TyJ4MHRME5uOcIejx
F+7lnetwUoBYFPzjAgD2SMLoBFrYsd/QSMT2A1Rbo071LfwzLP6MmHYvxDPG4diQylejD8x/elU9
P7o6s9mnlvcp6IEeXnwJvDYOoQq00MNu29Hp5If7MrWH6Qvyb+azrFjKREt7js3lZgg/7GGkxSLL
V9PR86Nq5Dg1g9sx5kH/2yxfB0qoogI8Bm33RfRk7qc6XjAQ/pV3+ICZ6tJfT2AOHhdXnJGF5hsd
fOiU65qUD9L3VQu1vpr4oRjRrGy6yLQE+Ra6WOhSMBu309k8C3zPe3HzQZcOPw/gHOYiMaEeBP5g
Fhz7ytOtRRrep3ymHMsHPxbmVKJcQf31UFO6TArdnkQAfPnSl++gBoVaAtejeFKn50uTZaITNt0j
DYFT4bXOxtdGvnQV/bmFpEjhH0iG3FWr4PpFPOVsvQayQcOldf+IwJxfii3lUd0LGYNShryLzidS
eePpAmUvJvvHq38eMzVWEVo22xpf77jO56xP4r4gjNRZ9+SmKV2EtD0DrbEnKeLT2TulC3IEUYiE
ES9g+wvaewvVyqQ3LaM+CZVAQ3sRHKZDX3QWLyA0UECk82N1EJqwUqX4Uw5NS4GKQ1FRbQB+eixc
+iYfVHEub7OXYvqoLSg8NygZd8a2ST4xyqL0DbKhIfGo10jES1p6a/eQ94pO0M+t00IAAiKyoCaA
Z62lsVN82udXEK9i0KUpTqSwSaeoo5wzB8sxCp1p0ibPIIifcrRkEgaeT/1deg4Fy6HkZuL4fP/L
rpVOzqCsaTe3+gBAf2/AlJgFaOC1zcAN0IIz2Hsl+noryqtF9WjOhBFAdks6x+J2IcNn6Oxgv8GS
W6Ls2C14/DBGelYIhGpLzy2qZWdfAbb+oj5bGQ2g++xUTYYRocAX+VsDBmMn+HW7Fw2ntMxiB58P
3z3hakE35JurYOIjmqYYHwAODJpxRoyYRDtuKUMAIKsF4dBrF1QdERCgMWFb3kq3hWvV5fhT+emt
1HYfaInDa3OVfLF9K75uou+w20KwfF0YgTc7cXYjJlUQHerc7Ypfwn+SRsiIpfafTi1b+/nKrBnQ
AfmTy0xsWrbNGGudpDsHDAM1soVxYswUz/gq2Ql7F4Mxy5w0+FDRDTkBwc4KDXiSAnKYLbVqq1XC
iTrKOpVwmlooH13GtUzfBZxZT0r6lWor00g3n0FSdxCzbK5X3HtzwFjyCZeFJrm2NVuKR2jHxF3H
WZejk88AvMwRM0YziRFxNsOM8djLu9f7hXNSuekcafr5Ydl59C9Dw1XKtjuVx1AnXCwxjSzg1Of/
SmY3oRPKcRN/kA0MQsMwfv1m+LK09b1w23bUd8bJ+7MddwVP5UWej8Pf+V1kbz++eMhNyZhIFZhv
KHXf5NjMQvc9uhpzYaI1AqDssJQsaLjbJCnZhssXFfYR+CS5uyTERnr2hFWHlLgQb7hon8fem7KF
aok5ocrw2QCLdvmnfzkzH4FdX6FqS2+utJtj+nrBpEGyQxVx//BVWd6FCcsTGX6r+Z/8pKcM6jC8
PWPe8hLIfZfm89fOuBkpkdsh+NfBrJfsly8OMusgukznNvFvqUzuT19jthHMb9mXeLVDXXV+Oyg4
1ccwWuv5TDA1NhHu9ty4Uxj0rW9lW9QNdO+UDEV8ayWIzSxaEfyO9g9vggiGgxC7B+15bXZ8tyQ7
a1CGQIbFxtVGmMQr8efA6G5ntJHRwMN2wnohDMp6gMmABfRNAjtlshyDhyijsQa6CjNuanKYo0Dc
eGJnXAWOiUnunRBapg2p6cPTGbKfcCu8PVMosn9dcqxBOjPLVTVL9mBx1VLYfWJ6YbWhB9lsAhN/
GQdFFNg3cvDh2eByRNPBv7McCgENTXHDSb+xXtfWuJUagU+FzLN/v7wrIjdD7I0CPF3M7+KverW5
FtKTHeqSMWPRpfxG0Z5Ws4BSFMVSRUhA+/2+A1no6amGL+fRbB5daRFrmlKEz87H9FI5NyIBCrD6
Yl39MWxJCXqbnGKj5AZ6tonat6yAlJhPhjIJ9o/jxs34Lc/d4NNwClbVqznTeSa4IRqtJZYQSXUB
pJ2/g95sDOGK2p6ZBsNH5t8Y3w9QT3AqQNaNA6A0j8UpHbB/dFZrk2h4rBtlhHu1YnBPZhWCZEbk
K78Zq0vd5QJeUNs2dKQKvmkfIqI9ZcbSUI3APEw7VMDpe7bHR1zOKLRUk3FDtRhCw5kX7Bn0uV5X
6rFadYUWCSg3EOerNvYlVRY/4sPjCdJc1GBJ4MIeKxEB8hT9DfbCIQHBAxmSL/HwRkeV2Y4Nnfr/
N/Zv4hQPssXnxcpqg1V0nc4W6ln7wzkUw2ft1ag+efggNgtYDWmUmwOa69+zNepKvJGDYo7p3OZO
4X9ezax7Zi49bw5S96+e3o6s7KkjzLCdQoByuDvr6KEwfVb+zfPN50y9fHFQTHcuWLFa25HmJFpc
si281nMv2gYe3eUYb7zbod49MB879qlQsHQDH7DNsISVYkgYYSGkq6X0DqtoPzXeyuCDN/wwxDsF
LbDH5gjyF9MWL17xt2kJhrGPLuLhnQ016O3jlMA3EToV614Ip6pr1+vtbgbomi3WzMiJ/iLOMMww
WNsjpmUVWeLBg7Sh8mJYYPOwKkpTvJUXpMmjWJaV//5B6LL7VNR60ACsuZB6Y8u5LATsWikn2gkm
QMAjXEkYkAluHYF7YFQqx9TC34MCVqfBHTjJ/vovc2LdGNTz/SupFv5I2zXzLoy/aQDNDNWQKacU
svvudlvYi5gkaQHJboPqNQvtsJxWWO99W19EZcKBgRQTDyFszd4DqtHIWoOWdwscIpdjPNnUJj61
Spu7ytdfyyxAiBBk5snhuVCUooJ1Ax+rATAk+ubrEbSFTugNXAoUlB4GSpsJBJs6jx3zmwUiEbS/
PW/Nvyt9JvMug7xrCEk24qUgr8zoP/IUwekIFlaZ9eBwFz/uudQ4I8ZFExB4SfYQbZduY+uCBSmh
bNjuxtcwx2O1U2z2jXSB0U7bRh5tSiypwVjgz7IOHe/qGGL9CYkeAahdMES2zNmqu0YEeHgyZOpd
KuQztN5Q6pxWKMefDFS8cEFgU7DqZtqLnFkm02jnVCV6WGawWzozhBC9n7oNxzv+ZmQxzFMR11qS
pQYk7ciKc0Qkq7iOmSxC3aYGZYCt0EoWbhNtFIocGNsmpbLUyUyRbQx3JLkFuWjVCp07Q9mCPpbf
wP0ubMR8J3f2qv2q439qRoyec2NELyvWnaOGjyAnltA6v4P/jqqxmtF8oiJXofAio8s+RlPQDuGo
5Nf9e83ceDsXNoNlyrsSxZfBBdMzcqJiQQiI58kxTiurDWbRS0ssZq3YmaMRwmqlbUbnC/Ckmht7
GW1TdYP7hanBd/YvQjGCazTFkGLd/mRt5mfb2668L/TcC2Vg9A/jTwfTs/T8DFSoRTwFRWXOM6Ao
HIP10InHVMobd0C3YG1tR2ZJYNhcgChcQqG2E/r1FUnklw741eqfKA3KLMSklAE4yynNbHpaffed
bYY5FgPLI8YRAIm0NPKk4TwFROLB6SGD/EiheOXCVjeISzbBlwFOIXjhedeOgdICtxcEzDzDqrs0
uXE3BLrAmIatzV7WrcLrFQHAcBLs1WHdvjnLnU8qC4gTkiD82gKrayoBduadiSYVlmunRNxxmOmx
09jbscWgOlRlgHgS3hq46g4sxFprzfVqy1EKq7rO2PiduxklcPnUo3Df/6wtlP33gaAuK8j9nTH8
orXzJS4lx6YUBdYO+85MVUw61Iqolnjt65Qjul4lTu3D+ZIpP1R+eya1vrC7zqNIFxG9klApmqG3
fu+nGH3hfDnvFDxGN8z07KUyepbZLIpQNFyTbzhtQ0nwnCOT/rIM7sRpBSKkFf00AKDf5iSSMH8P
9D7ZcvPYOVQ6KoNJK49EWQRp6vqyOJihb2f2/6UqaByTA9GPONbAuUtLV3dSqYfiC2vrTGTG0A10
44FQCx1RwDsETxEC6DllgfpUQ2n7KQimYsdOfk8LNZWCiZ/Mw/CMxcQs8ffxoP83opG2624niUD0
MaTxP0shvbskR7bEXclgdwNEgxo/maxqo9lTuDnA4zybrP8/1EcwRWY9nqYJd3ciF/Ll3xF93AwX
kcwvihxoOV9+WS5/RTioOa3dqjNpn5lWmmUIKujAM7Dv55IXF1AMZXpSDxciXDa9AXnBMoSPlQjk
nlbWjWurnIlgo4b7wkOCa2YPlukAqHkYsn9mACqoC+ZM5wpdaUlx5T2VhCkY75TrII5wafx4KLTM
wRbpIfdyOcfeVyM313/CVh5mf1Cn3OQfox7/CT2neV9kAozjHuiE/LKGnxg/IAyfxst7DAA7DWTF
HIKcN1E9EZQJyHDNv2xEDur/02/FjLNByrQb+AYrm3ow5dnNjQzHsfVHL8CRlw2pb6RKUrqCE5Wp
pQzHhEuEcz5C6GFjBLwwt52sUBrZRVNdk1uZFPa8L63FZjKwjn2g3ErFMd9RRFVk9mtvalz15LKQ
CJVJsfFKuaFcEFLIJfGD20rcDnyl0kk7/9RV4rKwmlBtOGr8gwo0AbkqFceXcJbiUUB3yKHj0FGC
yH/CkthoBXX7EWHlFZvfPCwxyl/IaFyjumLjhH0n4Tso2JrLzhjMwVXb6iY5bbmiDA4WErt2YQoj
TZGpeddin6bBYdzy2vqQezQGEtMCvOYmVLffnML5fn0OtUKdwMkhNcWyJ9VD0MleStNsXH9vqfMj
snm3WHLxQI+unPnqFynq+ryVwrxI8mRoW9DYByQVVZdCV/3WrvtVtq3q99lAY5jh1xHvwbrE7Ijx
9RSv1m4mRCpdPy3Wcyzb1bFNFkXg4FH+Q9Q1Y17f6xjgRrOo6PcUHYPSOtfSZOvN+qL1luHC54FT
/4INvAseyk4hoQcYE8tsZKMLCu1J8e55Gvxhk12QNkENKchF79RzSxRbbFVWCU/y6AweSl9fbS4Y
OBS6gBU/psX7js/HJSFl5f/6WZwKyeii5PyPh4P8xdvPCRl0yvAa5QVdyhF6miQM314ViyzP3YFu
uX5+O0nSM/JvY6iVl8IMCRjlENBgJlgYTky7aPK9RzerMl8UJTFPazGfbOScz4OAlCWZP2jinC4z
n5cxSVYUvDL4OaWW33JpWokbLx7BEzpejAv6ifqpIHv+65RIrcobbTBz90OSfO6ljfxYyJJwYx3N
0uU/4ytmSxBSfKQLNsjS29jFxUgaiNGkz1x4QW/LPIraDIETNaP4a7F8jPElxT8fz/8EXq/CcbUR
CsXvcajTfrniKEeLfQ30DwTmEid5pi0WiDZTC7AAVZdl1NfCIpv9zPOoTMVQwR3nafdgksPg7K2E
NmwHWy126P6Fhf7VmYNYeHiKNMrLFHHn/Mf02+x7t7hLZ18IQp3H79pExGeRTkegNvlIao6qxdiq
q5AEJxM8lnO4pdSg4vbzVJzmMFszHT6mXhDimTpuRblN4kfLr3IwstpOkUHwjHhhF7MHn96n41nJ
e9bIYkKD4zenXnWTwUrobiTdzYCy8oN1um8wdU9SWjo824VJUh3GD7Ynsj00qTHelRphFB6qzE3n
Os0DcR13wW19dC9Knx+b95lbt2A52vH17sx1zF1Gwq9KYeFZE8XRnxNYSelrYBOBXH16iTKxMyjX
yIEMQ+WK49co2Yspx9gXpxTDVhq6wD4qrVGQsp70gcmIC+irKvfuN2+kgx6+J9RNz3ms1eN+pQAR
nq9MkQym0WlXqHKZ9BYPwbdG5T7B3ulrHh0jTcqfleKOpXvOyHunWVVf5kwps07hs+wl5G9iPDKm
3FhjP/hoKB5i8Arfw3MbMkms7fzvebja2fBnVZnOkhchrdhXPz0nwkSJchbDT+VqFvKItY/eKAUy
jfnPjRv/CfWLoTdaZaVqSYgNr7qXXRsZgLXRkczoFwimcT2dMQWNzZqbXXLRQDdqPasCqkiLSXBw
fSlA5zp4ifGliWrL+g1YcO/gdCCOm5RWd/qRfvGEFXZGq7cGzx23lVxtNV0gm2C/jgOSNbVqZT7w
2oYeWBxgC8+Ij8AMcS0xY8I7qLVcGO2xWMJ7aXCe6Ev0BzzwYL4WNvc9/HhYRbjWbBB1crCFv6C7
MNKO6Q2c252WHY36c5gnKK19nnhnRVzZQ1CqpH3S6cyKSHEmkcQ/JrjtAayWydy9fzdVPF43rHf5
eix0ulMumpzNqH8nGlfjr8ZKAn1h2DUOZE1rFTsCOdwHTto+FpsG9ovcRrgHOD5x3SR1fb1KOMhE
oGhovkwn+dgW/luO3Ow+n7e8zk7YnKqmnctQ1Z2rwdYAtl9aYK4VgxSah1XPtiCgTQm9ZAEncT5O
K+wpAgcMxEvQIenV6O3bgYWjIbh3VnjnvUTxtguF7BIipX5sUJF2pJ9SheJZ+paVqQGGiya2PNfc
v4keH7Akv0M3fRk0QtBUS4gMavshlRxtasd7eonOsfiwyXKmcpj318UeqIHzAKyNNeAda4dXMrWu
2uCrFFo4mKc9r1it7kdbNp992VnVLFb+aIRb2sl6S+Ep6U/0y4qQLo/FBbiqutfzgvuxEAsFgsDJ
gpUyAcm145WVt0+PsZsncfQmOgG+k9PZK272ZTwRS/hw2/xe+kbrpLvGLqpcVDww6RQff1xbdWRr
vp9t5efGJyvAoB/7xyXwJDoIPKo3ug3SpZ7u1t7TbpP/Ds34fPshh5zxupXT+RJw5YUuWVu6565q
XNaKrXAu371Qy3gbHxVqZn0rN1KN9Vy3gWA8pKR1KLn5qnllZOSgNEb1G0YxPgdbtLYnAvcMU0R6
jonlwZSghqU6CzmhpwIhhsZf064aWV5jwbB2LJ6iYYeNPpzJDVR3LoN7Z8cq1w1abF5dbrYKlfd3
QMUOupWy2X+/xbVddGRGwRnCSnGJlnFXFVBZ9Jup9Cj6E+va1oZwnfqEEFPHl3l34rQEu0TVppYP
Z748Mb6C4zh8PBRy3HTk6psGlHKBPMCEQJHYbmLJxnF8p0ZIlyf45G28SZzFmzp7SFbTWI00Ho/r
rPlq7LfasQQUT4Yczd3JizEKMh6m6cx9X5SqrZQw/IveA8mDHp+Lm0C6oa4C7lCCTEgsC2tsvDvl
lDi3Jbal/b4Z9Wx/jr9WJ3vSNWKBtDDjt+bjpgv7stOnued6AhE0quYu11/Ob4667Uf+G4aonvM1
nHtAhgPT9HIb6lpVG5RQfqRGn0g+O7qkMR8w2cKCL/HL/E7ibebi/9ltN8UQJ3tAl/UXXSXqUDSV
Vn+vLepAlvkPZh3p4DuLocV4iCBcBAhz++X085FQ97nHmALCJpDdTLQaatSzYyGx6XldMPrwRCcK
wJN5PsGTZTKSWz0LkqEhc9no2FZUyRmrEKZ5XwDuAH3gTqYyHBpyCtrFtH8uI/QJYHnK78td+wQs
kdkk2He9XyeYQOzXlx0zmjMUGt5dDiocM8mAY8yFFSKNVt7xOxbSJdPUcUGAo2YZ0/AldhOhb8Gi
dzJMjpP66gjiNbjcevpGY+++HS4JNfQ9yPpbsHBVCAD/2NI4m1rm2LXZqawfNZwaxAXipGsT/4Ps
6WMrGFxigdRv0t7zJWeqf9Ma5SPrhsRbFNFiFz4cgdtWIRVI6iK1GGRgovhh4Mh7dMAjqGtdDmF7
pN1IJ8zuvay+iBn8NHgBH6P9c9/9rOxC0N4WmygCSuSYgnmFMKHtO0krXBbbZ+po2QTz3bbvt6KU
TXE3trzQ0g7efY8S7H/wrldc83yX2nY+rLi1XcHRr43uMD1TzM5VOQdugeLkL65KULphdyEsa+bl
BeHf369fUaOFgKzRkqHx12ULVAl+jLEZi4w7cRRM4EcC2SpJfU1N+ZHfmPRTd1pmIf4OU+T9Hfdb
GjLN5jJHEogiSBTBRzfGCWB0vAoc+hKQXR/6l3D1gKRkGhBe3Jrl5w1A8D2xOj4N2kR5l9GaBGjc
zhwF9h/Lq/4WtSIOJFSEaMKbd5fMOj1aobYma1A9XaWLv+HnZEc8LJTcOgVxQs5DsSXoLBi9ssvS
gSdF2UD162XrXDPFuQg9tXY5/BoPTpdCu+pqtH5MSeICCGbcpRqr72+TPZKTBNugG2Tg8W4QCk9o
TaTyTj0XqtCrthLH9eYioEkgJ4tcf9l3Cpzj8GlenGFmUiYOe5kjvTLZEUKTGUfHkE00E6gaZRz3
vFZ9B6go8L6uQs2rGPtJOsahhDamy3KwxHZybA+jyaDqR4X+mRO1w2ErAwXsM3we4OorhHE/UO+U
Iw7UsT3Vqsd+YaBMtMccUmuMTW+dUj8Dlb6a3XD263zGlEzujf5O7l+XTKhCwQu6CzwAQnVc3ati
gas3dmO1APOxfvQr9WEs9zzvPZonhOkdmH4yeR7EgLFsC9P/qtOWyIgrUxLFGNCKFsNJz1CLLrjD
VcVMKA1+htRTU6k5P9NKvLyWvTADbf4xIcFLMzFZeVETuHP6+dMEKP/SQsWBFEotR1fJxVyr3NGQ
kyqUsbsO3QJ10bcdN6/SC3D9opjMuHJE/YOmdKH4eU90IFxvH6fuKtlepPI8SWnMiOpFQtIswxvu
WwXyUd4UIkCNPnFqMK6qTfpfdjCT2U4W0iuLoJfLuF+TGGv9sE+iztBLlhj1dtPIU1LRPrl5YEJN
ye1X/xjLYSBWQD5viHG9GldxYwSrb2R4M8inKAJRlPN6ghi1MqHS/GzeY3EWuY5iibkFua3AzebS
2HXE//G5ZbO4tvOVlV9IkW83JWdBDHprRx4H+t6Zo5tpzGX6Kr8ixWE7wy9aKJ1Cx2BwHpyAO3NS
fRY9FnW9Dxo/cImKBDkshXjLB+vP76TPtlzjV4ocTN+YSPp6X/5oyXDpws+U/YqtLtapbCFGi6WM
W64zQyGJvjOvRdfkb5dTpdjLcu1oIK2HYQ2p2UKcMyIb4YliBvl+yJxX3/ciqDqB7pFwthOSzh6e
cOWB0aCuJBblpYLIAqwtdFsBthLRJuHo7G75UnoAV/JfK8zH2CTLu+1+NCtlvgyvpGNCvpMEJbD1
cdsrx/8xg9tekGnIMOhlgt+YNtSLy9yW26AhlIIYF3tzDvwOTv+otV3T8HRvXeCtPTGM1o2pJWq4
XEB34mPnaYmUklEM2kYFhH22Io1myIwUU0fdkGMmbS2QbIZ/yfMiBzhOLWjd+oIUljSvlY/x5bZV
D63aGR1kbtKEXZaTbYaEObIQu11e14BLt3R8CiPFxVz6/pqTWOQJ1VIr72r0OaW4qeJ3EPtE2UVV
FJcQdWQry3TyNGa79J0I6duotCZ6z2DqdpN8UmAmGOT96RtXTv08lyZOZ5STY0721lVyocb3dq85
eNvZmRZL79A8AtqJTf4u1UXAHmP2eJ+QnH6go0XLtI0v0T+ws5C6yBPYyd194K22m5jl1ukr/ngi
vY2O/D2L/LktkGEpMK0CgQO+Hs6efwYU9ytCTZ5BFLjpDPnfSuzx+K9biXqGP7nM/Y5d/RnenruV
uSncRl+idbxVtRIeRoM7QbMFaqNhxTBfaPKz6/X4vV9kHojHecXF3qkXFddTKu2bcN7etQhy+3vB
DCL8hw1NSrF2O+As1lCjfEPO1OIAG7xCgr+2SHzJSG2uNbbjmKAMxH4FL2+G+aLu967O/Wh2t6tY
yoWXnCXXGGNw4x1FLjYqmr0cHO66O3T0YqGWhMD6K3C8oEMLZzVhLogimE+joHhe+YqcYh/oEl51
YELNEfzBDohFzgxkfqWbnnKMiyXERHHSz7X6A2j77IIhrtDb9PgPAyL5Chs5XCIEMaHTUk894hn5
JVewEeHvxobZkT0OqfSvyUXPqNrXTTjXEhVeS4u9TbSoSCxahJ5EN/xsoDOUchTUK4QkoSi6Dl9Z
MkT95Cud1wEoQ1mMhr3Q0Vs9GKFXHwmk3h7+kbwvy9kEalv7CwjHF0fS1svMDpUKgraWwreHhy1F
oGMCH39VlkxmU1HN+ClNxUToaR3HpjfI0dL6+HfO0a9H8NSdg84tGN+Id9rBuA2j1Alaw9R1Jje8
+WQhsc73SNBV1eLP5SonvNu3FEbUoCKMbSyet4uu+swjQAQmiUuGjtL4n25nPNG5b+2YnMiKVBQE
RcTCPC39mfzL5y9YhPBvpD2MHdiL0G/RZGr53u5545Ho7XH/ki6L7mm3IHydhk+ZGVrqjNymBulv
h5V+U7yrRIsS7lHchmufQUrtKDqPgdr9Rxk7GbmWptN0Pv+dfhmcE2nslpnBrepL9tD4Dtr6/VM7
rKSqFKlTDm9FLzEoPdHc6IDwm8IiinPJQsLt6F926+G7k8pr7RSuMNeQYajGNzZ0h8n7WCKFkepP
1rq9Vkgk8ez95d8RRdwa7U1OojuZtwc4fG6REc2/5wi8NwJAoQdEqsK6lGsdO+RuI765r72wSIOh
Rmxtet37HXjeTRBDYfK/WMSLbZRiUzNFXad0m1l3Bmp4VYfsKaesWXgztSuE1kui+itiItGVbt+v
sK7bF2y++WOA/wOnG8JFt7u+j0sqtVTWFo8hZ7tp7Jk504g1eoiN6Imt6R09cfLwpF+fN9HIYjQC
EQrcRsAoLSqz4+mls1r8UyBDq5FOirPhxxJVvWS0/oTKyypKCHCRntfYMLo8uEC6Uba51lT+NRMF
j0m18b6i9EWAwK9VvVciPhR+rF1k9eMasIBse2sSzYmUZ4EV4DE/FcwvcaL1/6CJv5je78Mmqula
/FA3GbzL3UgLUQtft9RGtGmx77dokQj56J4gB3J22KwN0uccRCa6s3EoR/COV81VD4Io3IuR+kBk
txVCV+TCr5gAa+9tERYkmowkPRoh/OTh3CFyU/uFxLIc8AGVxjNkh7fjejNIwwUIV68bUi/VrVha
6qofZEcqZ9+bgnFPIqZJ/bVHiuF4Li+nrePyjIPlUxcpeQoh+Ta+4HrLlFZa9FKaIITe+L0zr8yC
Q/kTLPDfhOhN+TePIBqT6NXrbIm/wka6T5p2ef+2/syBayea0l4fLuj17BBTAXDkZ83jjN1WnxK9
qFn4rtxG3wygloU1FIFh0AsLVFjPLrVHbo9XZoXhZKhU27f1e52jfhFJTx5S21KgFttn0+jOfHk5
2IzKXyxoS0qEIr1UMDDOHNSyRRnVFHW90b+7EAyg8w41UVvVJ237FwZ8cyXkg1zHH6yPr89VUXCm
hR5sZAirJkWR+znJdnvcbBd9Z2f7Kvx3HAu6NEPxAySdxZiHSDw06iEhMtlbCv/SAKb7SpKaByKE
6AbibMN94QOAbc15AufejD1hVvNkthup6GRn6LkZBOxcVHmornvPhkUTNAp0JA92I1k1mIlmpAhZ
Zlzeh3pr2bkbuX+OrTKc8wxO4zCFuh9BRZNfhBmk55xTUWH/ojWnge3GkSGFIp8/0MqCFW8vaiwx
ozc2DLRlIZH7ztMfgj3T8NoAgG0wIGpLZfosCGIOYW6f9QsqxRNvA1XeyNb+CEJalyNebo2/fkUy
KNBGrmIJvlTFeo4JP4jtRNtwdkeKsNb3MGatHu8e6OXgVqIMQTjBPzxrB6BOgG4vfozH/GtfNda1
9t+12uxjwMCxaMZH6kRoX4tgBcnFwRAsWiUDg0h3HmlmjgAEAAB/eox6XCtaQSKMCukoHmF+TQ8g
1uiDrephCUQX2+CgdPwS0INvxtZ9PLnTLSOTBqL8xsp9Gv4ibqk+a5ZHgIeDhaZsuNALmoXtJRDz
zs8HEpCbcgI3Pl4BLG4PnRcmhNQEXoTG7CDaix5P4a1xBeE0nRTxowL2gHEaomDAZ+JZ0DIupOs8
c/oHmlnXc9QMnMW1nwBxZYViV7sV+z5yfTVQjBGovidAIQZiTy7F6HhdnFfw1zDJQ60Z2he3OEsh
3a61rmno5XhEcHMpKxNG6Bu7dZtIIig5hUUSyjcA8efGL7MNIX9nQ5NivRZOeY9S56c0k5Ennxat
4QM2qCVqPD/5OmSxdiRPpvSHsflCl6soq5pIQTaUqc1xNfj64rqyVroZRs3yDrU50va7DrI5/Jui
kHbx/jTuhlUrVdNFORG4pKnQfBZIV3eEGAYXoZecYzebsaqTFmQ9GCaXMuSfJLAx3q8OqisnEdC4
h5pAO6kwxnEwdBqF9t1znh/nSW1JljO4I3eKN6z0eylQSBZQBl6QiPjLx3D5eroq8YusOde3k6ef
Txw5Ig+qxKW3bD/HaW4T5OtDEemZ94mdEFddWYOzmoDQ0MZ7p0p9AyHLDkpta2dRiATpdyXV/IMA
1nEiZUX3lvzybWIJAJ3o0JGw176IhKhRJkTbnSbZ6HWd79hrSOdx5MAslD7Chofv1ek26SNk0H6z
c5agsaMnpufmgLmPtBusmDV0Tpp9whRyeYhTvY5E6UArY1r9sjlL8gHe6BRD87OGVSfYuIJ3zcsR
VZzA9w0dEFim1a9gNRGb3Y3AgaKITwA+bCirBx1Alha3wfqxvMMoGtudMAzV75AwfVoyDl+7M0fc
r4l1WD4Tn8qux+eW85zSX0IBvKF7CBMFNRKE4r3RCU/+yug7V+bWQHnFWAyf0LTMbWGtJbeYghT1
cIpgcZN+rsDacj8R8FoAF+QqyJHbgHphBBweC/7AWIV49UVWr/R2U1seMANWAuCMMVS9fLhm522b
T99fQ6i7ZTCLsiRRD5zQgEhuztKmyWduWE6dUJLpCHW4lkMl5cYMP3tDj3t/Px2jolCNM/0gub1g
5/J7LumD87EpSNgZngLzfTesdZk3kM/R4qzhaKJY56Ga6Y5lUqc7o1enNJKIyslEuK2h0BWqdh1I
34jndWHMjHDlb8+qScD2cHvIn731qU/2YXtWt1OMCCyTX/qbpHL1MetK1psceJJ5GsYsZpxefu+U
qWhVdA67ztn4/1xK22lQWdoaeI7exz6oUjTekX3SOlt00fQMfuA54qZVNRUz04sAWReyxUkP9459
R8UJedAWu5F3QlKIpumpEBPwQ3puOEx4Bjf2nwAzWTZfznrus5m0sgDxGMdu0U/Q5LWwioWBGo5G
GxVBaGHrMhFJz6XNYAcXsimAc3vKxakJDLbLB7DIfa97YvuG4/5uC2cKapsf4vP9/a8Ivn6Cxpon
wptOu3kHYfrs5lB6y1vr3M1AYqFQx720nAGdJq8/LnttGy7wHR+6SulNawzSgXCBjiew+87P3z7J
tAx66Vh5Gd9MHPZzyL6preaztdT8rFBAi0R0YCxrefQINFNL4eBSmZNtylQPSZvz5OI+fJFDfXwU
1nrN0K601SL9vpxSYA+r5QxGvdkAyBn9kaD3ACsc2mWDWXZV8tYB5LswPWPCOWWyxvBqNm8xszWa
wyNa+0bd31P6l/NP9LB53fo9bZ9e0ibtPd9IV3sgczD56jBCrqRljmQAMqQAS1IbqQpA6Sg/BhSO
6yJPq7UsNQdNEgYGBo608SW0rGZGarbZv1LayHbbDGIDDbOEjcyXHxc/MBj30zp7AZWrcd3dwL6o
vjaPhB4wbzVzE9XZ5uDxtKd4kHjSdEcGm8+iUog+6bv7pRLYgNTibn9+McSxiSPIKeJir6mASQNK
cAwpROz11mgnKtftqaAtK5LgL0pcoqdLScYL/bjRXP5RwGk3lawIs0XSsJdKCWAHrkS1O/hSzK+2
/baCXHktKpcO3QndZaUgnYF9huB0XSE8yMPUnxUp0vU5+eamE+5tZR8UXy6/COXpx86gGNAl8cu+
pb1YRk2YXyXXXQYY6CM7VyVd9vQUAslDxoZzUYd+tiVkkaG1i7o+0r9tSXmeudmSDPG/7Bt5gtY4
d9InlivDxwG2URGBMw33FeqQ/iqKJgT+8N2mS+gfBNMs0aSOLQiBvyq6KEK1Yl5fVYC5q+56P279
7LXvI1WgeNi6I9mz3M2Uc83mXtrmb5PrLOFp7ON7x3q0HcpQ6f9rtHqoiGdlBwcas2fbrAMFVb+L
d2a8ISLMbDy9byHoYmM/jPi8dXTK0B8TsR2yrcFtbpEnsGlP2cyk1Oh4W8YB0leCTofvKm6eQMGF
4SegXP+3fqM4vWZaW4k0J6sUAccVCiIx8euqgRZoPkB75FIyEsFOuqsNgHZujt0CCK9GH4H/raIK
2naqLUnMq6ALEFVSAlXvsQpWkcUiTWmuz81YJ6U7rWD1H6h2Y+xntc2qi1C1b2Gg98A1oHO3V9Gr
qfmMJEfQIBBKF7trkKqcLt6sUwUfPwtzB2oyoAaNZDT4dv6oAV59HiTNFqxumWg7ptOnS1KWO3KA
d0bRvFVeGIe6pU652TQEmYZPW61be3uV/ZSUsyoTXcNAdKGGOCYhSriXLikcZ3HiJyppjqyHqbtu
HdpFeDSEUSuxigiFYoZvdx3qwmtE7/iBMVxpgua6h6wgcKuKyUf5/RQsvYcdaLIepUeZ+D+ozGQK
5vT8aZ0IDHBblkPQTXCKlcuDQomb6wJsDpaVen7cpF1f8hWu8lM0gchTKj6mplhjCjA8aHB8ReP8
Poz6sLOzuaFW+I2lUfg7UcCtCaaiAhTvQ4LZi6VHKX9TkUWEa14SEgix5rdesERCz1TWL4/m07F/
GPzI86vpMV9rJ+Obmz0GOc4RbdBdDaBMNbZ2NXM3/xLfk4qXz8RcfBF6Hz/kbeYgJM0ntRvYfPyd
/VdcqDaPJd+bH7QGzyeY8ZmtQgWfxcw0ujkYHTPbDdE8dkYRxIye3SDnkW9wjtUXjCUXjfRMs6uL
CWfJZqQ15tRhKHmcOz4wecJ6sTaM6BtEzfsW5R2d+9xtaNAgr64vkclksYe9cbqQp3dxxj61g879
NR4XsSqXsFqSwwQLVLh7j7fRZ1U1SZP0v3Q8U52iwYS6jGw+IoUsmEAhs+G1WX82zcLICKxCHZ9E
3TLz1geOLYsysTed9eZYMueOlNhgLfT2zpsfNZc83jlQFreYgrKqKbEApuEnTyM6MlgGU9SvrSpD
mVQm0VgJNjmOTjezAubMd5sBbaPB9VX3e82C859NCi8v8z/XnxUoc8k4dfIXyZW6YQAcNz+ht+if
nNIugf22ToClxRaCRm2EAhyzdoHQ+0FyIoN2oW3IpGWiCNdnkd+wVuk01ub7pzUO0nd+4gIVzlvp
VMrRhwM+GKFYFjLaj/SgQrtPzjwby0AJrS1BngDiqRXADjV0H5CEn5onD1BBr8oYmFtX15rQr7Yi
1xFbllnl/QyNdj5QJfhFqIOy8em292SC1WGAOfSNSACDg5z+fx+T4a5jgGoB5HiPLDb3NE7rGnJF
d53JaZruoMlEoHlNAAEoIFrrPnoNYFURNg6IXuMdo6ldqsk2yEPAxS4tM0/VSciV7yoEg86BXJPH
1Xg9bWWCOfi/hHc2Nvbej/F02wuGTEF7qI1WHRjzTcRa/u01ByXGGpYIZFdk96FQ5vSCm3aT47uC
pMYLbqrZ20z9glKa4K5siB7ZEp3NmFnDsILs5iFKdNYu7VdG45M84w+rCToWzSHT0idvOypECy1g
ljE0qAg9cmU7vGDgRb8TOg1BLd0EjqdsJf+UuNtdCnq6VFf/eqwslNWzRYPx7orqftLrOJq4rG7K
JRtmipaxHnrjhXOfWldY7ZmKOteDEnDMc/LTScCXjEtBUpIiFS86wlUC3d+STSuVnux3R/tP3Czw
ogPx5vCVvsI9aDt3/tFajBiQuJy3hZI6PqPZLsN42W5eCcyl3DM0Pokl7jQEpad8XoBxgX9OQecg
Jvhv+/rIx+euvWz3wsG/Q+ls9f2HJG9ELPTW8Zz2SfE8kmn9LGjhDwQlAZdsT50jbF0h7QgviYfJ
ytJvcPOtnJV41ipg5GBGtr8glT4bVmdwKcuKJHmXcOd00i89/XrVI9vSvi+SCEWE8Tmzq5KGCOrp
kxvQW5TIhcHzwjZGPBg+SNEr1w8l5D/bKQX8RLjX/LW6n0mSN3iKMA/Vf+Vs27Rxr7/s4ABGGYvj
zSFEls9R96cBWRvgAC3dheyZrx6btBrU0o7J7sNhycfV+xBIx2L/BiEi5xTaPqt/Nx3FkXIDb9T6
mEi5HWhX87ZzQrs04rCWoBJ1D0sZ9R1QgqHbtHNTR+KLYdzYuz9Tbrl8P5VmgJ4CTcRyFK9tI2bn
A7qWfYk7XUyFj4CViseJUQJ467gbJ0fNgq8PjK3JeFULbsgot7BE0gxbvykpdkrnPH5EJ/FG26nP
svAKu9ot8uyKhGyq57PfuVyj5AI4KcR43JMALHr70LhCXR2L8amiCZVcZlKy1Ak5qdmd72tm2IoR
2mRtT+Iy6YP4GBwT2rA7VYTKcnNJ38QVnEjqt3hfXyvzJWuJ4Z9tcJPZyFB6TjI9EH9PJ+d9F/fr
JNpAbN5IOoxwpUZR3bGKHEpWnQk0eYvqBdvqINTl3qhE83x1kM03tXAPLjneUUr7glFFhRcNOuKR
DdHKMyC5SGiI2b4moo89YSl+eoAFLb5nnMdp+36VDP+WnHmHElVkkdoUt8uUe+nPLK2+GFj2id6v
rW23m4PSG51/Y3P9UbTFZ7xlPQEf7IfJmZQ49JIAigNqiOEVa9YsO3t0CsFmppTixe6h5G2cFNfj
V7aodP0ENlwLrbqWlAmiJLN8eI8hG/wVvU6z1eQk3o5h8sSmd2c6oxDJ98N587Ss0+ou7NKeAe/e
dLeBcCbdxQFvtDrlMZMCdBlpZua2FsH+WPSVPks6YCiMoQy6vR4PE2Ll8sm95wtpiicutkaEyBI5
7/DxKltjjlOj+SXbV6RxyalGzquB1V3gSoXh5p7sTN3r9fPU6W5K2z95TLj9vb3jBZqs8BctQs53
EIhqGhkgSOaJLJPAlq4/LKHQ7Y9PNQVWGo/Lszc0XflJWDIRXsQbHCJWVfudMnRnSVFtK8kxmHRw
8CcdaDkWFCyVzrIWS1qNXmEc3dmdhR/cNpAByQBjGOpzas8qnDPA6dzUYWhME1c/cJFLRiG+r1ID
mRVCuH8cDBJ74K5zoauEUP0gdoKdWUga1KiyKf7R2FsBaQOI859khUlLDu2mj4sOIR/8aOOXD+oT
tWVU5tjZ59iUzLY5RsKn4XZJ9zCLMVTivfcQiqOfGdY1tlAfmdHcC9+uQK4qCUPgYxywcliCqZ60
qYCDXfCIlH5nmj7GD7e5NreUuUSUCybGEXaoRevzAtuktdWZi4KRBojtwqdHkwXb6sQc1YMMHhtj
fIrXbpMzwlSYPJWWp7Q0qNRYQX06qdkyVE6gXLesdCR5MbyykEm5g2KCHqu1lA7miyn5JfpWrxvu
FyLQF1DNZmq4SsTZzjyZ/9SJiWhQ7wqqLNqRuPhX1L+cKyww8wzkGJzEw2/dGMfHVR4EwQFb3Vor
fQuMKx6Yon0EXtnOHOQupvShsszz356VKDaGYiflOu0Ws4AEs6Qr3t1C45wJQKsbAH9ihcL278Gg
xMXYEkesV8qhOM94/gAzUSj3Kh8wF/hid3YsUBgjyG/pNIuH5T27iD8cTstnroLOlMpYIoFzNdQl
StCdsQfWJf50VZ5+3rgmz2a9BryFsiyuWQCviKR+584FeqRaIr5C8rcKYt5yoBDR6UnpvEbzqlpT
zKTQJTpLhwAy0eHspe3J//4MBLZAuV1zdvW3cV0SZURH06W5SmXvXw/DViPjnQd4azqEg3AGO7pT
NB5lnDXnKd9PXfqmprXycBU0D+VcwMRkNo3fhon9hPj40M/6h/szy1K89bzFPcI3Kn6Bo9wSKrvz
kASYePZZuXGSoMYy8QYvH87PSC41C56C5yZ9J9e96iP1qwrEIghZsquKDuU7bAPt7xry+t1lk60B
eSImJ39tcGNJUDUEUB2XngIF3SOSEVIds/19vr7D8NVJ0siqhoUKnUfTsuL6IDl6bwQGRf0TzDS5
y9YhOUHHnzJom2dLpghjFOLB54Nqo6HOCKb8TPjIdpLv3YnzFpBIKluto8GXm/6yjVGG6ajXgJ1u
5WlbXdvQORHkEs2JpyXHNgWOxD2uKYqIx+YNfpGLCzO5ldQMehG4SoFxUbixggh4hMY5MgXr/YK7
uhbz72igFr2xxDDJG7FdSsA3c7WeUezk7dxzPs4kFKSyxVTO8kERnYf4N5Oq66ohBIo5MZ8X78pa
eIR4bZbHbvz3hAmyvS1qdruN+ZCvb4gd71OUsvJAoEdaHZJZ2pQbT6BdY+aq50CXaXZJiUsjw6PC
BF+0fRac57rFXfhh1YIQ08lRJJPjfKGQlO5bkh21+y22bQfKHbkkOCzse1iXYcUdfEaOv9qWTyo+
nHbAO7XXtg4RzWL04s//4afqFys5xArZkvqi/oQCxyHmZ6DDBqIifK/lY7kkwgPgHZMwfmm4ZINs
gZTOy/4+zDK+ElpLJR3saSYJ6F+Tvz7rTfUnKPP5JBuVhxppWbmKpG5h3dGq2PhxediHhyrSoXkt
DJhYhXyH5rw0/wjGNH++Pk2nNjkEXzBmDji1uBAstabZsbtgujgzZbYid93GicWpyK2OSUGL9uEk
jUKRZOlkxzrdkKeRCFCytFILMTie2VG72+GI5/pb0Hgv1JVft2+keluLz27tmsauXw2eUKKX8nNQ
wi1ialBel5FPwgecevh6VJFsdvDsnRKv+NYxc+BtEdp6vjva2oOWoXpFCH71xS7bwkak1YyTf80g
OyajS+oRmyV8/7GTZJdZQeVu41Zqtge6RQYRwi9XHyxs4Ysg0/u1nwfq2UIxSX7XTGZEWzMmI6o8
4ZnQfR8gUWOukfqBEWnxfoa6kLga1ncwy0G0sYuu9di6tZCYyAArfavGBMBtAN07ddn2n947Ym/K
iuqkHFQJuxATIHiiT1ry1rZNVKlUne5OSJLHKIGu/myNzAvXmElt4xVmrJClrx4GLQHCi2nEDSPr
tLI8y+A6b5dadDl1G2XcjKyAjwZt/iU7cFe6Lwm3r32FUtyTsA/T8XqpUeA+I6vqAK6FlctUcPaW
xQq34fV9T4oZzMef0mxzQ8oIwn2Yc9ybFLTkPp4jtHGagoGAG3hLaA4PYVPcmgJvAsvE6n+WSCYv
D6FM9A+X4aPMRrXUEb1mxvKYlqqdp0iM1Sig+Zl+QzoyvFyhIjdAccqbBsGn+rAdZE4MXbhcvSpv
8IWmEhr9zu1NTwyjPV+WGQZEQ8tq09Jf2yi1H9LkzpSKBOrybGgTw48AjxNLrhibO27Q6V+Hcwq2
d1AFc3g+2NSvnR6cY6Ejq6GZKVh7JNNUc7QMN+7evD6L006PnKa9vGmUmQWE5Xpcn3DWxXF4WBEq
2oPNq5IB9b1J2vn+D7a7QMT39DvtMl4e+MwzEVdDiFim8sIthh4SfDfdA8UnL2E6LH53YKZKeyBf
RlWlPdrArkfsg+5NZSU2J99E7LA7u/xtGF7oVJl0kf5y8Gr3D+WSbmQrsA73DHVtj9Q2ENt+t0BX
csudBDBglXf4232TsajutnMebo4q53ce33FR3NzF5YSdWZagQYmpVKvkILnPwqub9rLwGCTVilwa
B5GI85VCkFIc4yovTxfWSr4+Owj+Uf5A0amZ+FzC3Sp0ofbMYS084OWHDfVMOAPvE0LG6w1PeMGz
WWsHpQVlFfYk4qyFBsTsIbsoacOnET8FzF+/RlqUGdg3nV+wPT+TJeuIig0JasI6poVLhjbh4Dol
Rdl8q9ewExyC7JJq0Caur+CAICZPT2kWexvftci95UAA6c5FeRl64HCKSSImzgJNFwNxJIesojmx
FSyf6mMxSKN1R1Dc4D61BpNOJ0BehiJMORY8dCscDtHMdh+nSnITJUrl06be10Sa+h8X+/1S7X6Z
7Kx1sYpqtN4FOBXXDpz4m5BpwganrIEV/8NoNK29iag/Fhhl8ioE5LuNG1VfnW8SXwhvJsa6TXkN
dcd3pPlmmMr5tdBa18PR3f0/CBQoYrFu4oHEm5QjEbZ8WqNSgfQocwEfNi1roa0EhkKgF4RjtDa+
CMRjJXWAy30RripYyj75nsINLo1RFY50MRlyxwsNvMGdClwWE7HNru5Fu7HQWleqwzeyZrCc81D5
9XsToi+G61S4PJ4W/1aL4cHhoAUT/pELjrsnfN8AlQ/ai3/5nsH0V1sfefXHyQ9j34IfASPwhoJw
22oU7V9DlH4581lSzcRf7HpSc2bc/9SBULvZZAb3OJU/pjimyChDiq85xxiJ8bXJOQS2mUlOp468
ZrdO1K9HDgzziscV4A36aOpdx9or9HNytekn6kmsVhDqflpoQlmbY13yxXJbuCEXEfwaGR2ypYhd
SV+qgjSqdbEVnEJN5ovGQsMB8HyvJZ2UK/jIvBnjJnGqddm0tF+CqaP48PJQA7E2cOwz67xBKxuE
6riT2bScFtHSJs9l6TU8qePKXOvnMCNwrWg7h1tRyOj35/hDbggmKxrtRgZ1ifxmIHR0HPSwgiLI
amVZj2GjG8eBthKT+9TGsu2zpTyjOGbVRnFz1AEV0O+AMDjklwpxf6HffPP+8qsFaweR+ZdkcGG1
l2YIoI1wWKLSPgXOsvwztLw/ymjxLtGqoOGZAvRZNWpjIRQYH3/uQIZdZDYFFRXzQSyx9Web/Z3y
lGt1c2C8lqy+5z0Fu5E0pSAuLHyf95NNsy0UnHBEE1NNSEiJBveOybeSMB5zA2LIdUjnNyK1rOUI
1O1PPa512YvWKXFapJAOD0MZtIO27raZMq5jracVr71eL9/nniBEPN+jEvnLqqsI7ooYWCzohSwG
6LRIC9wycudBoi1oFOAMcXKG5E4e4W88bPJxh1WNvHN3bZEGd2IkkpkXZxlZIkZVEmsCtXQiZvUV
OhUiOxn7HRzG8opDsGEQ6XroE8nt5RQv0NjLefx/k+7S9tC1IJUajY9szNF8cpeBNn7wLaeJBAYW
IUgTjxHfoQZcBKlUZAZZgRK0Go8kQArFbqRHNMlOL6hIuzqtKm13YRb3e5utYwVTWlB2zz/poR1T
wC+/IIrdg1ZikshlbNd2kx7dWFeh+uqOtdeZD2ziScLnByXQ2fb0APujhU49b10RTmaezFdxIvyL
fArQcH7NtQ+URSDBcRi40za9KvHNXBrJgzfvaf19M66yMVnaI0wKsBBFsVM/vN7hTSKATWNaFH/j
SjF5wSW4NysKbijRuL+jOPAChz48pCdRNPl7G8+nFREEaXUGiVPQMWDZfvBxjfMgATwfcdZzUNIO
lQyc+jphYX59jOPHfbz5BymnonoPtMG/XagUcR7JkS1LLO3IJKJwFOE4KsbMijjbYYsRTYY5kkF4
maFt0SWMqbFp2rQbBUB4spbtipSIqcDalxZKS1FPbvukM+YsV6wtv7R0XXsCkVPs/Dzy2wIDfhq8
9zolt5trTDSgdPQy4/jwscZoNBX6gnSBfCzdddLyEdV2Y6zmVcBvysZ3nLo8vOET+oMq8jvF944z
GKK9p9e8bdJ40gZHo7wf9mAqxBsk9JcblDKGGrG1Jm0cGk1NzRjGH7rpSZH5MPzlJccxKiMRZj0O
xsWuo0TXzCmWvOP6XKel1jOrKraikv/LhLOLwyCwsVxlLznLRWKzA7wgs1BlKoBgXSEPq+OI46/z
VgqmoRMcege6sxdNWiT5FbFyXhEkzDO730elrQb/t5IXVNEunGh8tZhKQS9xvQDw2xVzZSkUximU
Hd2wc6vSOY0OKoSNUZqjt5ERWHE07LXIHRkGKWhUnCmuPzxeJS+4aUJYGvPPMLt3xuv6YwJRmYqd
dWlpbfoI04FHdGceW9gBMrIjP7IVa/lLcFAlrLkYUoprzSJ1CYhKLVztS7lRUKfK10w7doAPWtW9
1NEQL9P/DVFMhrsIyxUKCLQ5KkGBlwkRDqbewAWhWqTtDQEHwKIZkqDt9n99Ah8aHDmhH4XjrHN4
g2sW7IRTOT0xvLYHrhJxUGJaujXxcXeFtQ0Qii8zumllQ+1RM4EZ1ZZzpA4NKzXGtMVr7TjWaNXz
yuEL1HkOoD121r6T9ewaxwZCZ77evEhjQ14D+tUBkSbGwNEwMJ1giImW0/NxnYgatXG1qmNSoNNt
LoFOo70hujmYVBKHavEuICHgsWxWs8eILox5Cj6IvHCnA6i3IdKphfozWdk6q0Q/POfbfiN2PlG/
9a7aaKgiOK9bB2kaU8JRm9pHukUx+UX3aEQhKnPUV42mMvIPCJmizcDbaEFJU8WqhAiPqVgWrRRo
bi51mZ6CzzLlMNamEVoohDi/XrJg6SUN4BB3t5RPiOv9irRbw8KIPHOUxEl5iLzkj6vdvdzaBMFA
/ipQeL5mpdFWpRaZ+hp9V44bgPjQ0RgjoUKP6KJmnuZwtopXhqZcDlB7X01A46iJQIZyDvsVkqR6
yssfAnRkpxEulAtJvTSVSHPwL4MHyut+utq2lgI4w9jjqWd3Q9f+11AUUFVHmr1GrdXsVOiV3r/J
UHgOmUEYCbTug0loLLIiRDGfnMqEXPZFp495iU3hXu+nLWCbY8FPfzhoXpJ/2rNO2WJ4DxW1v2NI
2gtygg3cgH62UYeQYfM6E6mBzgsSsQYONpFs0dSuUo0NjxAVQU7uiuM6/216uzXXec9bZ4/QEUPq
3uAcCURemINtOoHSNtL1Z3m9LF5CJZvh6hZ+5TGmmtncTUg4WKKGIcfayJvhiMUJFqpoI1TSAfOM
rtIa0ZFJb91QTMAr3G0e3IhQ3yISmejnZ3TTj60hHnq+Y2SN+YaRFDRwrs/zlA9w+h5bZ43yRTKC
L8ZMvUAtRUf1goHl99OT05m2aJAvUryLlAJemJXsYa9pfhfmi193dBwhVkMwjlOozajUPiaMeGBn
P7wcLhuKw8f3bmH8bICFx3zGhE/8r6lLjreyrWjbZx/mzmwenfvidplTMUgO/mAnYD0NMuKNh07F
va+IIDUJpwz1OScPSCVBXspzjf9S77eaO8DxB8K65NYLVcNg1oLxTC7eL/0UelaUJg5GBb82Eqpm
sqvzAGRhVfmxSSnsiNAaJR40v+lt1HcsjWTEljHDqeyn5sy2wmT8k787p5iAPEeCTqXieBiN/sl9
tZwvLkSBShHWwzArPwr+peig2Nb1mmge4e7Ugc4+Emp87EHt6E7ugfSjMPYBVbWR7WxuTvGDr365
PhQDhJ0HtzM+pqP+2WE6iYV5Lk91xryVjcBb8cF4lf6irpslgImm2mUxrV7Meqy6ju9mEjIccNzQ
VzhO547A57Z/R5wibY9b6/wFh2eeIQniyCTk+yu5YLciUhuKCv2tX/YbzGRklFVSU04m9mjVBfdd
UhbpP/PetK2wrcBYfJ4bd9IVrBeCWOBZ3dpDr6BzO5wfBzpgFUerZHHbza/X3SEpyRY3NncBoxJl
xtDnvUjVt0CEEpSVm7piudezcAFS3owSr8EdqjnAnlNxPoWHyZAJaY4VOxV5u7CwP9jIVgmRswN8
gKgMzm1W0XPrAfryHjczCWsNcvDEuCiEMJ1OpAMYv20obj+by2Dy9LVlxauASgWPYW0ejf2asgxn
ixRg0EDELIBlLV/fFYiEpd18+zDG/PSzNYdC6xnCExAXNjCUQNuKZ2LZFJVkzWlDKIQBRwoU79/8
N6F88Q1Li7r734DT0paysS49PQuqLusMbQjl0Adjsue8P2k55zsyN+PeQmORePpglLIXDRcgNLjC
qkdIgDFOp+RnUm/NM6I5T8s8SQKoSqUm1rWma1IGq97GU6Po8zj4g6QGjL6jp2vtBUuLNwfcI5JE
RAHCxyUGev0N+wKZyV/UKn9RnYpG5BhW6pAY+A40Dlz/mj735FBT7bAx7tUoLPfg33zBXXAK+4/2
axOutXv+1gEAuRLPWppaHkRG2XV0Yea5NoGVjij21htpoobQMFUxMIITTaro5nsO0eKF5j3IwsZ1
UTOofovfv7HHF0DZc6Kvk6E2+o3kc5QxUUKeyLI60eL2/6j5MUcA2eg4W562JyllR0OkbqIISj0H
oC3rVkgeyzA5ya9kT4IQFc1z7nl1sz1PSpPOir/oxMFV0cMOTB1mgXGzWub/r1NoTcazYsOoZujy
IifGG9wh/36YNfackhc+hys2Wt8328EecRKi/fCN7Yav+o6WVGIP6RkIdij5wTLkc/bEgd1HGUnF
h4uLd5+U+JRDfhkZAgKOOY3hLoBOHFto+pAGQMZWO9Ky+p+M11SWqQ3USwORHuPM06t4m2rZ6OCl
BqnMZcy3jM+GNzdBlTTikz05Krv2sVXXFyZtjrddSlJswTlzUdZ7MZgVvkDLgf4SCxq97kxT59d3
Ai5d5dZHffBrJFlbfQBBPPq7EvHLqq7X0NHpRzp/51KVKbzzy8S1xd/eXUQuT1fQwUH+AhL/eAUh
QlebKW1BZmC698B0mj1pN8ysEhXeRvKwbDi6IUc0wc1cwCSS9HAiNn2C8g/wNuoow4dMH/hy5I/l
qsTaoZnJ8TKqiWA1xc+DCvFL1MKvFnDbF+euQFSxfk/H2BXdBPX8KRN03tJ6oqXcUHcbMaxaorBq
sch8xQIaVJ90ayxUGcc5MoOB91kfrypMobfsb234/I6a6u3a3qCL1bVqtJABl5j1YfJxbuX/93jb
BkfFGEn3vshV+5pjDKJo7ARARAmJauPzo9IRw5CodwXSJWVc/h2dkMXgUsUCYWplQXi+wZKGagvD
YqJOVszxlDuBOXJfzC57o9PSgifcXprDjxa3kARGWCczTfhO46i+z+6QK2aliXP2xRKuOKsXEqw0
G2ltZpBBic6YnUTt6yOmew+W5YmwV2pOT79/aOQBuV10OmqqPEQHIN2SIqOINUflGoWMaKJ97gI0
8euCKTrLQbuomOho7PfS1ZuwYRtfpLwph3CZmatRgt32kSiRDU+OjALLoqC5arD6PdHqNfD4mnnm
2RSntsx2DximOvjGaJczqV/fMzmuy29hRMWP+ETN+cQbLRXIed8b15E62HMFxqQmDjloVzEHC5T5
6+jgJ/pUH8MV0+yQJD5rTK3H6P0YG3afB4OFHTTy4prUO436MI8ADRCUXsxwLO6QGGWKsq/jRomF
dlE1EXQ6WYuE2c5Z3Be3zd0eSjG78nomR1jAYUlLKZHIbv1+85IQ+nPYrSP+VuYdUmDyFf/xv2Ra
tDjK+Ay5VHN1vib9vFqubrY5bYN4T/cr4F+W7If/3sORxPw6+uuk4hkNqGv0/CzJRzNjbFCT4Uvo
pbNn+yBcBZ38STSW9Ftm8m1c4z0ils+07QF/zElufU6Q7vEDl15MQxQBOPAKli+EbBgAUzWLf9EP
fT7eqwwpj0IgQEMr3EPlYinGfiRP07jEDEtxgV1cym/TuZXXRvpLGvtonKGhb9YoSouifjlxPGwU
0iYFbXMDRehv1OAgGdGkfzRoOI8VB9eIogyNpS9rzKfjpWSpZXD3PIZeFHBHi6ASehrtz1d+PYe2
DJYGJ7Yr6tGDgFz0MfKj+wpMMkMykYSmfG+IeJpsCiCOZOyUshcJ9oLmHpmHRw87LZPjZ29GHIvx
sR+HUqM1h5Q5vtfYMvPCn2LwR2beWQZdmB7ch/WRQs0zOuPm6n2av8gd32IVnOW10tnhBMWgXgjF
6prZRBkaFGH9m6JX9nBkEF2to+pORw9ySF/oWCDzrhxsMcUFaiVp4Uzl7gMM8r/PFd0dvPS3vBU/
e8NKEGO9XGEYFrsxuqbeWbLkwK/+AqBPLj8jPNY4SNXVekVJBbWtgUtyN6hhn/SlS1tNqPEDPPnD
6Z6YVMtZNL2XKsoXnjY4u2GLfXq7jRvQ7igOQPcD6MKlCXXicUXcd7Patu/o60ZzZv7riW3ZS4zE
bqiArXN4sKoqsp7byJ1mdSCpSeIhsm6gxsxJx0DmKQ1nRQfx9B+/M7yWvB3HwvIUZX63xhe72WZU
aIa7c/ivr0eomlz4goY7cupQ3ThYBPkpijDf/1fERWwfwz35huUS7TnuQ72O6QQk2jSifkazQo/+
x9gDrcvOUiCEUOh5yHnc1P3EXn6QhAxRtQ65sNmki48ZxvCYDN7ahK5KrnLT9aeBuO6B1BoN8Sdy
PyLREpxuff/8rpS8yQAKfxv2cvCYxQ8oYepmQPl73ps9kDKM4BqnV4RD9itEtOo+m0Plalub3KFx
4gJ/e0ezqa7ynCdvP5UR3VzsauwGDzIBYPmPoVT8276Q7MRyAAKHb/pv62EvPAuYl+r76xHs4zE9
zJj325S0LtF8JGPL5mDvBIk/zjW4rO1g8WwjUG7JZGj24Pxpx2Mthg8YDFB697Vf2cUP8ZLmFAMV
YmydbCwNPkZ+F0tWu971njBbUG/KNwIFkwwTu5p3Q21d/LwpseWCaYeAK3ndh/CXK1ax095PqMsI
fFhoHH3GLWiXc5RadKPe+pgT94Y4cDAefSXXmrq3kpADUQepjJBbt7xoxEdQaEGLt51IbDvn/348
ga+poVnyfsGpgK9+kQw0a5buDjxQPiQFdxALne9l87F987J2NiSqPHm4qOz34J8nUVBXLAxyYE90
LizhQCVLm0UfyC/82qnanp+j1WpCr1nvC8Bsof30lPU1VSgCDk+VtdwagtOXXMTVUKUxLRTyM5H0
QfzWWG/FYdcy9TtwapNwDZvRnZ3GlsdKxW8Pg7OZiVWea/OuNizSwEb7NpEl+l1wyiryWTEgCpsy
s8xxHowlKRCPf1DbHiHHzbEiHKXKhZ6Jw6fQjFNj+qI616EyCT3Oa0g2UoLI7YlWtcoaOvkIYIP3
85+jD0EN7znkSmJCbC6HX+Lr0ZR00Xd1aM0IQqESOkOR8nk7/Ml86D5eqU+Yd5oCM0bC4UusYh5l
PZ30aGNGAGcJFYXJlnQe2iazQv+ZuTvDFME6Ymkgd77h8NKx8wBn9pNxhllWxqn/Q74QzKDk65AT
okOWfK7hVTCQbJpx4yqZig+CUHo23H7QLO0vF/bLpczHBQ+I5Wx6nr4T3ZLsM3D5XPpGZA92rUf0
U5lN/+562FB+NVGWTfRLM79AA4Y8iZCPDhmF/8BOBHklXEzTDRS1V4ri0d187kctpeCCXQgeJ0iq
h21kg/91TTTWuuWA7bpkPJjUJBBnDmn12/ecJ3NGB5pm8XnocNXZr4+v+oZE78Ea0kMfPi7BX2cS
hvEBesb6lICq8D6Uj8QnilcsYeeM0cnwRMePv+YVEucaFA8/p+hvGNoIItNQTWtS5eG4aqlYpcf8
dDDJAoyEgLkLPS/2wYIxwK2ZLOKkTjaiqd4SEzqlPN+JvrOu/uKRyXWZpxRroT0L28CnxgLIJpsu
+4dm3Yzlxm3qXC7XuXmXmgd1pml06XYNB1UwrcRhaNURPGs4OLmvoaU7+Sswu6Oujs3yMhcEXu8K
qoMNWngbo5lLcWdzvYUeYksJChnzIT09veMhqHGPsc71Hbd3bPNLBJYTkHOujsQ6OMIeZTCSpsT2
e/XvoG+NxZkTF4tx2QSxoaDY3yOFkQrrT1N5eu9L5I3l6OAZivWIvE0Y+Z4TwtDNi4fKQMGlcRzP
u6R1IwzDUigWEPEami4m8oz5iLD7D/gM2Lo7p5qdZpohBajBfhiwcjCNpclHL/iGXIqh94hvBKA5
AsjqN+MbvHdhTTL0/Hgi8fn+rwlZFsX4IuRkYBJHTZwASo4k/e0ZhVXn/wuR8BqWwSZXAp0kpi0h
sBgrimAbf5l5FDfcBxn7gTGki5S04NtT80YtCzifr+Apxno/07Q9if9BwqCaUSkwWxyEV/zGh3tL
bgiK0+EUXLDbIZt6E3oovRK7o3UvAV4TPZRGpJuBVnnP3qdkcqwQgTopDbzqvsNqhzB2RDX5oFZj
YL110Jk59u9ijrIQNSIPu6xZ2ViEp2ecraqdo4qlZUCv2iAgVb+jdmb1lRxtLBc+MnYvqBjHFRx7
1V/9CTNgrn4FgQhf/ABv3qb5sYgXJ3ds2IGCLK0ZVQP8NrMeiW9fsu8p28c+be7uW2AV3pxQJx1L
oeNPooPK0VkoT4S6TSQ3bJn45rZdEPs94s55OnIxalrg7tSI5DjOG5Nl38bxb8/hhg/MuWJNyRiQ
rP9PFz85hSBO70uMM6uPX3ZVjpI3ToplBCFuiCl+PsaCK1fJQR4OXYURVuIXGviyx2B3/9FUstqC
XDaCKY4YKvUBabes8Wx0KYW45RSO+123uwtlZpj63qhYa0jK9iDbjUuEM+gtUm0eUG1TaAYEzFmp
udzj+DevIvAF2LF0CNSr5bIgVkvkiYkZI3pfcqWsHzzfEhG40R6iMs7leaEJxU5hnpsuAdXmF1p4
oj6iUI3FaZNTf+rT+1lBVW7Sz0Lz/ZUCkpZRfkEk8Qb/9L1XDyg+ULtnd3bKm5I4tguc9wJhBtiG
n3yLu8mrSBny/MVaH0VdvxAzghGC9tPY+M6C2kciZvP5r2CtQbZ3WaDGZF7tf4zorJ/+F/Tpqbj9
053jha95FK6P3Jw90Jn22iVVM+vxxDespZ+/tnWlpxyZpl3+bSsZN2gUUet/ftlgZ35Oe2Gh7uw3
gQqnxVGvemAmLZIAzBg8yaWqkttusoTY6Oc8rxJ4sIF/5QL+jMBCkpC/rxVpZ/5+wYgNujOJSP3i
ajxTkIQtto5pXrzbRWrVFF0UHoaLtFLFoMMpZQC+tbmvTmIhtzz8qJsviYB+UJ+36LTvUzZDuczQ
qmybhADuaIUC4+yRUeInws/yM1BuP3MGYVRxUjudVDw/jp8FMCTT3MXYWYo+YYX54utH7lMa6F6P
PdgacLkeG7xYT6x+QiTvpTnyYejgfWAwUe4AFQrFTyPz6sbcsTVZL4XmPwly7hlc5Q22HA/9NFkO
M9ec9vRA5nP0aSATcQD2OHIFRxMXicygRI5h9ODDfuM7xonusjEahHgd5p/SqYxzWBwbQ7a6EHvJ
SeGvSSIa5oUuiXyn6sdVaHTZ7NWZh1obprt9WB0clb9wAHZtMqF8DxE92x1MpbCWM9djd1Qa8Yq6
qs33P5US8DAnXccCjLIIt8zsrd2PIQUmUg3np+k4WboL0od3VPFZR1Iqlm+LOKbzqPVjVbM3sX4C
mYJ3bLJaycJZrRrAIII2dev2GLxJB5EJnSsXndmnfvIdMTp2OhYGbdaLoiC+iCZmJwAtTOL1seHQ
YGzA2wUABgmiRiR4GmjzgnxY+aZLhiFaKYfE28IkR3zEwunTL2zq9WH4VFVdoa8JYLJVtCzjTT4Y
nO1KaYGNYTLC7ydF4luFcNYnZ9jo0I6QhlC7LDVVrCOi7P4iyoZja96ouv5W6MHQZbNzlWoXbA2G
P7wDsE0djpFpYoIE1110BT7JUGqrMWtPzPb7oDziRoQ+vOCokVYy6+ruDB3VMmjYqRf2CAuZkAN1
U4g1vr6zoBa5wsebwlMF6WkUYPFwbfWpexK7HSlyhkhbnJdMHp9r4FT9i2kjEu99XpF22BhkHttK
TiBII8DMmMH0cJEykQk6G80QRwlxqWsi939hfZ10/8EPYefl35W/Mb2a/RcnXk2ITnsBr+qj9tkb
+ggu4Q1R4v6q30y/lTGF1Xa+W+SysiIaWFHc6kzytsPVr6CXerJmI/nr79bB8/kZY88I9z22k4jD
V1/nwwudeT9kXJTGvoD8RI+dJmtD8ofhcQV0gcZwdsjTHRYBDK3i0MaEkmHj9MTh2rI6aj87KQ3s
3ntxkguXVZwVyzYhM6JKvVKSxIdX3dHgro+yXXupLKs9smeWQtESpGHtIaXhBmNkPO53r0ygrfTo
Vq13bncbDEnkYfWtY1tsNQrMjzMky+TTlMrmKSL3BmsmgI8Tx2qtAvyFIRNVGu/qAOEyWtOzIJBP
mFrU6dxsN9RDUQC662HieZyICsb53itmVhPiEtWom8H9bjYSKgGRVWL3yLBiY/QBGVAqe0cYkRuR
vh9JM56fPN4fHuw2VNOvE8tXBQbYieKkCwaswyBBNMD2ADnniWLXkO6tVexPYQjf/zFktbzE7fk8
IakVcC+7p/R6OQ7aq0frcG+lRbYfn/W/ll9y7WvC+HWDXmAWJMbGtCQY/DG5+NRB8c6W/smGb0CJ
VrK+JWevMN0gjUvK34epnBOTtxu3nX2UTg/g9YKtgktpEhglOkeYpwlosc8+b0bPZinHs/93xMwk
aKzzmO7Vrg3nzAK5bkLPDYvGkqaUGpoo/f1QxgIlNNRUysda2adwlWMno/bJsfc3pB5mn9cs5xyX
G57mNEHLeaqPTyBnT0tmB3txbeBXgCzc0iiPT6sp5mQQLzO9OQoUjvkvdq0Th7ls6ZPKjqwhiOvI
VT4+TwvzqTtye7dlyW2B1sIBOYkTh+Fil65wfrZrjw5rKuGm87cvOiWbP/6dBQW71SgTFqRtnU4b
RWVe/E88HwA5N8be29urhWq+icW4Qg3LVVD0QRfhenG5XsRRDvmuiF/XA1MegxCPvwR7i9ek1qnu
uXa5+b12OTWAlIVDLSEXvTqYeoD5ZV9ssfs0B6n+1VSe24M2IRW6EK/PPLC/seU3Y7JMNKmsnZu2
gDnJk3KgdKOTrjxQwhiJYQ0aTuDNk8ReykUga1HufxFmHB2W5RvsIB8w0MrGWvYZ5SBXQ1RAd3sp
tiW0un3jPxwnYAZs9AHl2YkxXji5L4IUouw2tS0T7tgkDZY3SIKg0bnFSsjQAx92RG/9tGkBLAlS
KQ7ZYTj0qMbg4V2qtxElUxbsOjnSFjkJwEdcNHiknOeiYNKOYscDEix0L43LCs8WXhI6UUqA933L
ft/K19h9LDWKUZ6aHO1CUWtW60KjLJ5egP7+Hrn83AKfq7aphNtcr182V10DN+fjyhNLd58sff90
wCpsQpMgcujbhDbsfXVUqZZE9mSveSMBtA0OguB2i8mSp8nUoNL1LhNki0aNET1L9DhugSGvsHP2
DOiwPm3WLuvupvIi5b87/vwPqjeKYaYr/EyQ52A/s+m1l6Gz/Mnxh7mk68txW/ziCbN8k4AokTmK
2JTAeCpdeen48UumgsB1E0pLwWB18i5Iz7JJSmPpx2TbfmdD24JrSJnWele5WShXI1RSOxQscfex
S65r4KsZ8HPh7i8dy9wprmOXGjb3bTWOvMbl+Rszuexqop/G3V1nA3Oc0yD92QGSMJLAy/YlJsAU
3cLFGoVAxvgTlhXqYKicItb0cIz7dN2HkCPFUKQ6uJhkWqzGKwRfK15GK63BtISjHBn/43muCm2t
EMBCCIHEvMaSZ3T+V8Mt3aerr1M85T4JEalwPoU8G2pFIWCaovGO3wHMGuLFfh/xVvwZBIMYImJF
z/rDerAWBYjS51wMK3tuzy/KAEPknc0AtFoaU3Vy1QyntovsILRjTjxhhWS2RVldVwPWrRAxs3G4
dBjn1K2vcmJuMA/15JaTf2JVFjfF4KJtPwifYoeX3pPip79Lhprcq3qAvnkvuLY+o0VpSIOFkB+5
VYwo3oilMPBqJV+Uvh9E1zGTDPnMymWAsNYz+TgnK4EOfszcsvkl9XaUqL1Zx5/B5Sbb3otjibDo
Xfu9L07XQoCHxzv9GqnkamkSUaTXWuZ49I+VRR3ekNifdLTqxLMWPrzCWZZekHB1TtT27nP0R3AM
5AtZ87MCCFk4QEFSp2+U4yctUVmSRDLK+glF/6rP57c+XY79lK2cqERwIIQNdIYsw6eYUypboD1d
A05nZUDfa0aeL0Xcb+dLmrXLviO9w2dgKMd2dQhXQvBQ2AlWWtoMoVl9r6m5Afqav2XknG2ad5Kv
CCgYwgtgIc+LXoQYZZZk3tPXeAvhIn8mEd1CeiTc/TB1DDi26HDy1ppulzUFVnLl7SNArb4k9c6N
88Cyzg+DENBPeEifx57X4EmDXnar0GZY96ynPXwADDniT/2QiMxlxFZZ/v8RJ81dToy+POEpFveu
3gyhi2rRjZM2zggWyhuUZGV6kKOsM4AdH6/NsnLaRxnHwJkjBKT35XlHf7jBpPBqz71yuLgkSEW8
7vwd2rUPqFClxVYPesrHAf8i0Oijig6xSvR8i2oL1k5doFUKso+ygQZxADuSenxgeprI6kxN5nM9
4GT4wM6WSjSku8UxzgSwvZBXd9v3Vx8JkqFSX/UklaJlj38Ps1XZc/gj/YElGX9+ye1qFXPuq7Gt
HUXvz9ZyxXegY/8S/OS0QcTn+bXDZUZgrz47X5jO/MxaOJQkwHx0SPVVYlkRBc8qT7qTeJJA/2MA
u3qhAuk8ybD8W1xUifdyodzt8dQ54YcU3xO/9VofRKa5Zf0Pi2ZNOm79Knd7XxFwjtPum7cVY5wU
ROlE7ymsg4ZssjY0TEQSavofod5lsiDWm2hUjSssMgI7F7V+AgyyaKH1I8GByWRHsmu9QMyKTf6z
ZNLuaNu45gmshmlwD1zI3o3Nmkmw0Ktl4gLSvno//PuVnuhu6RtwfJvHmVXWIfrlEl9fHOIDUY3H
PiHZ+F+QRZrAFu3RehqRwAi5E81eHTG02zh0+MeSdThQJQqRTNVvfFSioUgMFn/1uHUgHgLFtJXW
7lrrMcn0GLwmoJazD4XpPLp9A8Y1OwzmAdpUD8qcvJfvSOzYzVSZEn9UTPW51ZwSmfeAiz9Q3FuD
S1NWd0v4Nu9PMPcyjUDqODBmhpmh17xfh83Ma3gtDIh34iJcti0582p86c/qWYCwRzG2OxNYFyrd
IbLBJT++v98Y8eSA1KbfnzUzfV4SoqaAMRMXnPD30fk4CwDwZeAsOG9BfzIqpS/hPCzjk+Lurtje
DnKl5pYcXJMV41FS3zmqKsGNuXapFeMm2jHyEcGdx/fbnqe5XtzGRa6KZcqY94517wobI6cyem7O
Glh1Qyc/FHafPCr83wZAbb3srkAYjpHl9NgIco21+sx85EYjbW+F4nv5OAgQwXwMY1um0jIAjp4y
G5l1k6Xds92BigklWubAmRHQpoRYJ0IOT1trMSXDaOuaK4N4hcCE/Qgtt775RFe8mubEYuwgWJUN
XrIb+a1E3Qc+/mECaQ22vhZY23qH/GLi7g6i3cyVWNHkzYzDUN6myCIIxUZS5y+tuselmgz4uYYY
pVB5nykpeB8BHsXjtGj/5DU84YqpOS4BsKJUvP6LRNCRg2GJeG7Q8ZgvhCHhGlUQMT1R+KrL8xE9
jJ4vKb+rmTRSitych8JBO+wXSnKpG++frCMl9hKIx8DgrjfTUSo57Xy4Ti3mpocNLG+E68jjA1OE
kc3TIAQ4F1Nm7SjyzttEaT9NjOoAmB52p67qVAknQfvlGTBBQhBviAFWg51tJhGu0YKYxAcq5Px9
TEQUjoyGTAwVbWs+lYFqRhlI60mvQjvKo1t+bovjYdI/gUX+65XSMIjlBs85MTD8UncxvyYHGF1+
eRrbjJcPAw0forC5s/Sl5QBYN3/I8y8iAaafcvdCjfb4hxXAJS36P5ygcq1jG395iD7Tvbqvqe2E
1ameZLdEoKM+LQyQE38/vZ8t7l9EpmveTZiA11Au1OcgL47UsSNzr4yO8rTVU9zsuuuFA98IC7j+
mmQba9FHGomg8i0H+eIqdm/CcsXB1iYkGkctbI67Be49IYSfL9l761qMHDRAErj6YiSIM2c1+jqO
PqIKd750myjo1stbSKkqJZr1IJrb7pcChxGfTpo6W6cg3RHFcFeTAjz5RGQL3R53rwFfIyFLT3Ow
Lu3FiJ4kRdfNRWH2S+2nV3ZY4Rk4OACOhth67YgqCca2bIF2mH/W2XPCTbp4SI94M4YCwA8fxMpE
E3TlURkarcPGk/lYrap33896vQYSIAzk2ROwRqw+SUQJvSGmyV7PvupduIa7PR2RvRpbnoI61zp2
m883iUm0u3LR52LlcR9NvBihKUbmGOOgCpuU4ftAiF5ME7aeRi0uDpsiUB9oYdgWW4LjI/q/RSQH
BuopOY/Jxj7HxPDSr8G1Bd2xTF/lcn2vI8p2vWjQceQO+7PYry9fcq9AKYsGV49pEd9Lnykwxcse
pSk1TOBRnYdKOI4IJR5SokkybyE1MRb4YbBvCOAid8TqxzpvRejkhbwW4xE548aaBxAxvneOOBOD
Fa/kAKwpFyMZGzNOSloApQPksBLtUW11NySUUwLXYoe0VL9LwQE9zGAeVQ1sYaaUCJ6akIP2o76q
S0x4vOW0zHXZG8WYdTVyzrhh3nCADHlBJ931X/d5ryWgLYf6C0AfPg7q9/g3UqNvvEjNMUZXdVzq
b/r9PC/lb9aJYJCeoaxD9Tn/uhiwjfhtnzOCkopsSTdU+UmaxTlM2MX6pq1CmGCJ0Bkdtwi3pjgk
AnXvF0aSiqEUTScwjThRxmiL8BTvVA5c19TpbNOGtXEIK2M2pub+GIskEZRUChNoPDLKc8piHFdE
Kx/+0L40px2GI/gybiWMwA6aEe79Qn75mgE5HYnpBvgGpmyB/LU2718jrnmCb+Ii9uEKhVhEkLlX
8T4JTZLve/UMn6GOgUmWmzWtL5zxXAUGft5vvVr9XFwUE2ZQQqye7XU5ilertuoMBznstU41KtJz
phQDdgUrwbveSGDoNi+Mh1mgLkC2D09QtN8eWypD1uzC/ANee4lKYcg96EdI14s/qcyPatl/vEM2
PmiXAoVxhqqYHI4LO/KSu7AB/MomEnIdBuNENQrmy7ZtmR1VyZfwtRch1yu922YTce+k/L6jQ/kS
ssfwUFDnuVhb6bwsReZlsIP/By8nTUHCrXzQT6W2OcR+HFDTWQmKHc4FfrZP9F5qhEdwoIvxpEt0
4Zieejv6lyeRBL/YoyJ2QIZ5oktHsEUx/eUWl5rOJsied9divDy2Yz0Mxw6DqHQSDwqoApLi3RGl
2Scrs9bXBV8vOHfpo8HJrlcnF0c5Ym7oHuJYsVipoAL09iFmCvlyviwqdqXZ2g3AClU+V0Lvnxa9
aR7H2oTP3Y4HW9t2wj4WCuH8tj/KD3ytE8ptEdr820W1PesQGALGYaBLQa8IBX1CFB8l/PmC+S0+
njpgnUOf0QkCqswjGSXYXa37S2IOH50SLXjMgd+abAu1CZNLD9rl6Pv7Icq7O8AapfsbbM28Y1Bc
YDArWCduR2jAWgg36cVVoUHdTiySjVexBHnbtf24965JJNtXgzCsNZTtIzjsjWYMa9ttSeaeZcrJ
Ov6Zg2SQBEB9/f2fGTLF+LsoSYc/wnmwy3oNfVML0zqF9KUW5BzShKsR2yvhoWE2BmoxbAgo9YKT
LBKNvZMvwd3k/uy58ylpgz8hkiOEs5d2WgcTMWIMv65T2mXyvkqXT/G2DJQlLpBgcfWrFZow5mNq
+T5XGo5LnmR9KiTo+dnWfqnjwozvcuH7gLL5ldft9O8Lm314x6kEUd2Gr2yUKiyKnWGQG4iAfZiy
SC/Y+9pBYnx3OsV21O0xXTvw6N8UKtQtgaSHrGOmmCh8+ZjpVF3dI7iCLI/omkC/cst+9yCoGZdf
lAm+dc/DG4WvAeJvtaxmUPYTQSH8uzbk+48H8952gDatoHuYVqhxRovBsz6b/Bb69T2BZK982tkR
pnckot+cfemI1ikZaPfGEiR5vpvR//nqhI4z3QenA1VIV7DIJIHSz0eB+yu3Jh31nszdIzE6AWzV
cD3Sni67hF9e4yKlKSmJbtgnCh8X4LCpNvvtUFOV+JlrwBr2upf2qeYgoBJmGT6SFsD5Y40O+rap
6beJeQZPIs3SGIuR+tDXFSUVw+m/O53kIw371AriYi9QIGPXclWCzRMzU+Uy2HpgSFnxgRBeXsOd
FHmZh4smHsJDsmIyZor1fiq80CGWwLVcY2VdrCEqG4n8ixlio+oZvtIbF0f64Nw306w3CibF4NdP
tW66opNyLHn4921JMjRbGfT88UbBtzx8O1+OVWDmrfCUSxjl+Gqs81g6EScJebjTxmhhDAuKH0ZV
cKEpL0sRGPh1wlh+giMh3n30AkxLJ/XyHbys7sFIXjpFUKXEuovyocaDjm2ijiPzZItUjSljfh+7
vOLYvbMo8i/gwBE49j01m7lhwAsvHY9bR1mpGCAWi7xeqP0DFE0W/hyTbBxhf29OKQAcsXb4stBE
z4CWBTb/yPfLKv158W+pUOVuKWEyET7cru8czLI0r/oNXnGJ+FwIIOlMcSATOhWnqqrJZCnorREe
L4++TA4vYckeWooHFlyJe3owzYhZBprBm2hMH68fqntY+tbh1k36RJlQjdaEs/iCJS+tYu3tNoIC
Jwi2XR97lhrgIAjrV9XTAw55nSHI6LpySJjn5HhMHxw3TSoJ6xPjCBoWp6DLrrJYAPfxANKJ++U1
2izpbW8Rf00/LY4AZmBGTePY2qNoEVtVXQyS83OZxx81mO6/MPNAV5ymBUJI6vdLmEOY6Blc6qmJ
1L5ip318Q2dnQFu2P/qSGFjA/NOKn5D0zVUmGhrMk8BYFPvj//hntbJBpkkGKyZvM+A7uGDUArZo
9PDDXVE6HaaZePYHdxPB1feokzSu0ceaGYXPB5I+WF92ZscZp2eP6Q0OgfKRqdlRFWrKrvYtZP7Z
m7mE/reyeK1AVudC6s7wH7UaJZaMvcXaNQjiGq151r39ZnPn3lwZseJu87rFe01n3mDPOqC2UHEQ
As2VCgh8uVusTJiJ7xJmhDuk4Iw2/PZgTy0btsFlMIX5yDXg7wP7/5f8NGGQnRkxpe5ca21oOLx+
SVqejx36w36PzvLv6drBa+eAgqtLuiMdiBkasfMzw6p3OKcnvxB44S+8dt7VAXAzTYV9mO4X1T7i
Y7ChrRLaQmrPlpE2AX6WhYUVYK3lnXwOhjBZ2mK/vOWirUicqsENyPI7eoU/51fgGzITuUI1X9Ig
YGSVJe2I6hzjkFn4QdJIjKz37hPmVBG4kb4QDegNxsPbQVkzEJm6MOKGMfUUE5iN/K1uljbKfF5B
MmRMutTS4hkjTOOXApHP5WGyKyQXcmjd5YnSZDxsNw2MEsdlz/DNe0NObKCibcN6bqukJcDDe97A
QT/JcVMiIuC4QXWcjAaPlTImPoA0XPHgS1+Rh2n1QN1pvc/DEOf9LwY5i9o1aZF3ciHbMhicYoqh
Ex7t8iWcFiA34wQh4rF558QDRY4uVst+Gfp92G/b/FoOSXPNfBmI1NDGL3JNz8aM/scN6zD5lIWx
i1lTx1gECP27aR/99zu4rOTr4/JfeJUtnHj/k6SdRydq/Okzt2S3wmCEJHlILlH5LbaUo7F/6aEf
Vt29YTS6ZrI/J7l+d0FUqAxeKBE/P1Ja9e7hVlyKuIpajFijDebpwXCreT2cf2q+8zrL1Ie72OKQ
2m94+UXlgf6ZpNOJZt5ZBS4/buSxHZdSUi2deb2bYJy+OPR22H+F2ZIQkRBHZ/grRachLqrjq/tr
Ihn0YyRXAMSN6FYL+RlOoGcqQ5eLViNWx7FBt8th3vk4ypnyoNdnS2V+mlX01ZePym/aLagZWQtl
9fMnqnWg/L90blG7P58FOqNnPCmxv6eC0iK/LsU/H5dwsyKTvYcKwiqPBon1somIepvfH0LyxfgH
FcCOjv7Q3tJDawJccmv6anVKnJkl0ub9mUYU3Zr3VLcB1ZWM4NhUx/791c2VIjj+IdORbzx4sYW4
sp6FJA+8bNUPGqkCp8fJL3clVdXaJgiwpJAIMY+1xNVW5ISiiCadOH3ULJzzwxp4E142SyWlUPQ/
LmyxfjW0BxlWQllPi+sBuCk2Tdx1bMGtLVFhUfZCf7khop3e1uq9S00X+V4pjScLpOHAr715mMMf
QnpS5dqBd1MTRVGK7Ot+WZdnthNrEgUiAU09D6rfBfRM3ZlaZ/tuWvqLbM7XC+XvBFnhbklxnWHB
GxbbwJmJonbpRJq/2nAOoh116V2OgkHNEpM1lfij3yXdgDuA2ANSeMuAHPXYl6N8yJtvjSbhEnrq
KQtBM1eDpTLQRShctSbugythjTIACo/Rx+NSXsgnbYedkTM/yn4AFKoHunWQq9zok3VN9b2skAWP
XHx1g4u2Kw/AwHqRxeeJdn05PtZOga5+F1h+n5BaUYTrVUBqBLyEFXJOSCxt/30mvXpqjRObF7p2
pYkH1faXY9/1KOG2+uF92VGNf5D1dI0mBcfXOeqe0fMrtB9SssOgNfbe/Rq8sq5LNQUcKOrSBvoR
7WW3l2CIqxSOAIgFCBBLfop8dhNJvLwg9f3QqwOW+BRHD1l6LshlH4oM3d8hGK5UA8cX9N34LUOB
GMSW8RQQCiV93l+wZs0JytITJLtiJwctZtdv2fSAksR/DSk/eFOCNaHBzLmnpRDhAKHd5I239Xij
Lhyk6eaXthx+g0k6kmD0+43AyVkiV454pcIPShqjm1vmRgU/xw1+chOBQJIv66MVWYyclqSszSrb
GFfHp4b5nv8RavgWOgjZaAak0BxQz9kjJfiLRE+LM0usq59DnlIvCwCatWH+mBjalguebYCazuCZ
kZe8elJlKCy0euxSVTRCsmxpNOq6nq/SVcTjQiKcvUUe0TVfXwetRJhXCT7NGsnq3gRUWl6MWQvh
yLiFwxDdVzZ6iR4VwQpvY7rgSHnsbQaeR2SuWYAjRnYv1GjHjjnC7sAuc8Z6sVpWVJtEB1roOVWt
rOpsdRHJEYQXCbAz2PJEBw312EoM6XG+sXfrgf2pyv8pBOg98piHu/t+g3tmZD4nNBGDpYA/PeZm
+RHpf7zuxYBIlORjgplfSVAj8NPIm4iQFM52s6+zqTI7nfgB41FW6Wz1xCj7cCJ1iwLBaH4fAmbe
dJmx0NkKUvolRPOLZUyECrWLN50noD2BiODj11PMdcRmG4zjBBnaSS2lxugxHt+nSChj5WVJtT4N
b9+GKat6ZP85SnjHby/BxOt8Y0BKMQys3+Dsp9qoS25JOczJHrh6IF6a0HDaJk1qNEeG9B8iq8dB
0rIt5cQ8++o17uQBsOhdynBRpysisTTDn+pBDqGmZGB29Y5gI8LvOc7C8/5q61cp+TbvoKf3259i
Pp4BkZuREz/bJDwT8nAyNFIKXMsFGbfDt350qVoppqx9DadPHi7AAL2zEu7FEcLqYX5twJsM7SID
sx5e4XqHoj5lamLs+QAlyfxRykHUT9MeLq0waxxD7MXieSkE71T+FZp1IWQiRRzBtXx0DSkEu4Cd
+xr8L+yFhx+c6cG6im4hEVVwBQuZ4mKpk8PUg+1fxRTPPQ5nUwSBEs6g9jxfiIWuSrIkfbxy6FkK
KocdOJAp/j2RKc2XztiXd6x5Tzxs81KmoVjBzOvuw105S5p/32Xa/cWYTMu8qi9EfLI4QMOKVqDu
3as5StXxv10F9BcnFteTx1XGYDgCV07mYkgaWxl/i2N/wGepehKGHZmbVXNVJP6f5DBng3yyxjMv
yQRphR9bJMy8Xnx9ELPPOvke615wM2nh1Jo6cZkfmSFtfLa0xzSTa0YyTMvUCmg5uzvb8kIOiMxB
Xe+8r7haC6ZuOgruTEkjrSIaPC+Dr9/o3YUNc63CARXsE/hcKDqX9hP+gqAL4U9e04s1Ka/CYAES
63SL7Rb+OgHRkKExepyeqiRasjkIiwVxldq3JqRb8hZnKIHnEXkXO3FZS2j+ypVSh5AsK/Fk2iro
Yle2BjDxCXHu9acbX5HscjdhDOrNEKibJyaSOIQMGZkwrjMiLi2wnsYRe7ktx2+D7OqzszbarRvD
NHEsKgNklT5It1MHGRPEss8vI9re1HQ0d3jcb1rGJR9GtB/47iIw0O5G5Jxzh1pfAKbopewiXXpY
RnXs2YBFE8H3gU2LoojPNMEJvJfbAJJLtqn+w6nm33NI8XF5kWCaTo2AVV8BGs/pVGWk/u4438Ls
LaU+LcJid3iYqYqq0keEQyLfrxmDtGhFtPsNW9SxfTsS+XLSoULBFc30+jquXq5l0VAx7aGP2pCI
q6dZtpe6BFZ3H2DbtRFl62trosJ4oEdWcPqd6rGP3mVDlfYwVZBdZzoAGQL6fJMNRV/ivuI8ey9N
JPYTOE5PDdckg2Par2zUiEBnVaKcorDLoWEd405nbNwEPHg8aMgOyUUf0FtwqF4OyKmuPJOu6z6V
FjfJG0PSEtepe5HzyV36+XKC5Rkc1qcfzOewx6eejH8NsE3LG0i+6iTvhUPgwbWyS2jpEIcZPQp8
IU4HbUVLNmez9tbMZRxwnFxnAnF7ECHOBrwcL71zuqetybhW6xeADs8+o8ls4m5cLTIlziOipk8m
JWUfjHd9h8SIlwwh+tkVvjP3wAy0V6l4VGugftD07WUzJ1+D22CIBlKEd8xOxNfP7i2yAVWHoKmX
zLPMR8qbGSh1GyYnnASxUebsc6sOuNYbwZrTmYYFkaWvMzHwwRJbjgPvaq2mPl+SHegRQW27RlYJ
UedctpSwyRm7vArHHtC3SCT2sg8gteNGcQN0yuWRUESviIe+tor3xpEw2vIjllrkZItmmdQMTQsm
qehpNxXA8hOvkNZUe0KQkt6EqLtKxE1bVMc/EIa9nHFhilj/E4+XLrhS3xDFbKa+9Vu76yYrI9LE
HYOyFIAjOm8nx0SmTAXlz9Fi6xWF0QtmnsSIgChDPHLvPWfiOuYAtZhDi+RXh8kPJOhTBYYNyhln
/ZzzDyEYkuFsL0cvsYWNK9zxUJ5xUGs6jNDm4KVbSe2h1cfTlDWTuayAm+51JOQWB6ASy6o6zfDh
PqjJ5KjEzcqJe1C9GjiaJP/zdc5MOBHRdENI+v5UeAqnSJqHdrghQu8FvELPXXPIvDoSscRrR9p+
7LuVVIT+be3VecdTjoAVGK+IPGmnaSBtHLWU7nrG07QEIPuX4fsqF2sNrbUrlZgi6+EaRSHlyYoP
WH9wNwVH3vVIN4DSsFLzDkKizxjISzVbEDce6IqbtFBFs9667vyOBwHWRO4MKtiO71ivMewcQ70y
prZKAFPJTR1pZqd3CNGTtkim558cWPaG8XSPmn/BsMwXdHcwFfXlG0vUEm5dSSqR6Bptuysm5fsd
ETOHyIiK9xb0d844dvDsxzimx0O5PYMKWkMFyFN+L/fWjaFgfwFhrmHSfK6lElHkC7OW5NxZcq1b
SoQI+hlH+/IIQwi85CRC/NpQuYOzX49VxRIhsOH6EuseTpoAFaSAGn4si3YPewNs4qUHtpFBZXAO
XgW+m9Kj2IhICJ8RIY2IiK8IO7QmFmX0lNFe4fr4py+S5GyhMuV1uj532G+PrPgAnL31IBU/0Bpl
zFqFhrNKZx1jdeXSHOiwFqfMJSkp2Z0/qPDz0c+ARCNGcE7iZGwP4SxJQFubrRtbFlc3Defy+V1h
dKO1CDpRky6SmxUGgL8/vdlEc+7baCgLvCjeY+/UhZRngnfCWCvZUMlwdhGaYyhl5mzNJxp6Ls7S
/4HTfhRa7LPZozGinF5e8U5mFwmqFockI6UITzb3fz+jO4GYLyr4hcrPQNGR2hi4RSyFx5lAMWip
hRDXsznw33noVBwceXRC+/DhZqMA0+PgUtAUba4bTopxEdBN08o0Nh/V9MWolLpY5edNmu/DpEO4
ihq8L2IrAtSvWHBIxQXlEI4hWX6EwK5qKK/uuX/jsizq7BIjH+fJyqGf+QQsWBsy86dlJKAtGJkn
KBrYnSd9O1+N1ZQDfXkqDse4d8YHqnHJ0zqGEoPScw5JPIN463oxLnro3fZa/Oy4daa5p3lk9S7Q
YO9887u6c2zXUq7gVhyG2M+8TJ8Psk/hei3KjSLijUqospSKYa956A5/khLWcIvd6AD9YNsjtP6W
4X8aD98IVTl78ZiVh1jCOm3Qb48XCOdzP9XWVRtIp2tEXjUqFfIAFmC1An1ZRDiMGM+dUqymwOm2
ob+75clMNSJCMqM0PtbevVWBF9szz16iM8+WkftEb0H9FyGpth5nlUogMToQzEC5uvsOGM2YV+cv
qjPaJyCf9Oo6OxxA+sAr2wcunmBgWt06rtec2ii9X5ENhLRPHQbC9sy2VBrpPP781nfhWnsngq9T
dIv8Zq5B0Nw+ul2zl3cVcdAQqHKLvW35Dt8qQVFPO65NBbvkuHe9m2i0YiMVASZvfhEDKE1kS4Yw
3tXdUOIJDnHDEh+VVHoKy/PCjmX11lm3VBApCb3+b7ya2gJ7RVX2cnjezDCig4nX9yi4cdzl/3fd
Hz02lfA7Oat0GTVvZvANygRS5BX7jkJvWn/eTjZ6LmHoQGIZ5cySQiEOleYSy+AxHFU6JOzbXWr5
pYFQcf3C6LDQPDVVSXIU/9S9Z6j1TZ7ObN94A7lrAkF0hOiNpBDSoYb6EPXyo4TxFNG4i6MXut5b
eH0AgfFBIt2pTEOreCtAsprirarHhUikKL3RdHquszNEccYgcMZZ9+/a1JaQLUnL8DtAzOVDhfRN
/mn9QKs1zMudzKuaxwZiwCDdu8APQVsXq50v4mVzNEvgpfiD3FMiPSH1wpa1kggoxk8hKgYDKqNB
CaAYgBMeQzHqtAvrXdKO54wdbxDNBjM9aov+o5EPfZtgHeRgHHLhxvMaVf0A+UzgpdH0Vum4AH1f
aUb9tz9nu1BA4M3tC8EnYNsIyaA6YgVDaH50s/Dh3TYd39h3raa9Lsr97gAddIm/8FxrTruHpuqu
mVafIr36gMz5QGEbh0DBvkBmDMuQvjr0gDkGocX4yk9lWhZI7U6pQ0gI5rYIV5Yq4ovTBgss7Jha
w2kMsB+CXLqL+gVPUlgV+nn+rM6YAKa3cdoDcGYZbtJLrpXj/flZ7GMB2FS4U/7dWMLTz+xZqWRm
yHJliIXqWCf0AeAmWjPipJOtifH4/WWy4sjhGIZe4tF2NxQFo7lK6f7cNoOBIe+jUHhTxz8TkCx9
8wqMtX50NXwxenPqOkj9EjujAUOoSYidDffaAuwpBZrs07D8n8qinnpfkCf5AKpv7e/0c2N39XM+
tUT/slvZXl5YrvEKdpWTAVt+80yVVUCU//W8cNB/nfUn9RzZriQ212JcwnKHMHNsPcvRjMF9kXbS
474awntCrQ091pS1LyupdtrCmICGlIY6+sZuVgSIU5Vy1JQGxN/pjpb3iCWeoXhXU1bC6MsAqfqv
QhcqJfGsMzw2ayhIaiOKe8iYbWqoMmD35Fr79xjcvI+7oagZRGkPfdt7J8+aWyyaVMz1WBcpJ1kO
KZhStw0i940yP1R6Jw3z+gaJVXJtrrVUSY8+JSD21HYGn1MJn6vhOAMzQzgddDnbXiQCZtDHtMYa
PB12zuJgcbi1GdNvjnvnSK3fSTzqCrCEf2szxmKz0dzPgMr7bCQHM+DZbehbB901vS+61Gv7e83G
euPF32cuqQ8y6XSlhACEpNWS/T7At/LNaEbCqomRW+5Wgy/jI/1pzjypegpcqwdimNzkNeLdwgBf
4qSxYkge3ZXmZld2LxpyIHEVRPP0iy5rki+/azoiEWhtNH30/TsMHpekiF+4Olmq6wSPaQzK/MNe
/KdSWrP8wv6VSL0m60QJDqPtQBbAA60Cz2Bqyq+MF3HwN6Z7bH86syyCrvRY8H1HgbUBoOQaWI7o
uJIdzNBWSD6jOiucVuxR4q5akcYWZIgU/UevBkUEEfC/cmTADDHUe0JvI+iohICC1Mdb6WU8GZYB
50WNwrhEuuDCQRaiuT6pjte41S9JUwa+MsoJwiGelP9huYv2N0QEh9jK4UbyKr4+SEzREyRbToVk
KgExVmPZIdFrZriYBLRwOF3fzCHCK7BjpNrWNu6/lfjGFwtj3r/R8F5q1s4QrkL2kfR6xqRp13WD
M44LSpf8KJC+Kcs57Jfhw5bSY7QgnNhhejjtlzVASa2Vow+8lgud7qHy1t8UGUkNCUrYkm2ehd+u
d0lsq9VyJVRwhfWuSz9vksfmxDJGBwPIvxSpVw2mBsAirZ3QhhBx+8jTbt+nY5JECSyfndWDS2mL
u1UEW7MTsEE/eo0iQjlXpvPQWqVar0/KkJbPJnY6A4StWVMK6iX2l+2iIg3TUPLtbwOrFJ5kHCqQ
LAnNWwmt/wdxhsg1PBpxH1ZRaUHStlmZ1eJFjAPOADnT2bH2Mu1TAZ3XRD2CpWdaiFt9iBFFhLWE
JLQLf9yX2vlzFMgR8TliW6qgpPi9pS1lLCQZ85G0QPnT61QKPmGlJ6Jr/RTDvu91v+BWVLgMlOZb
a+LEKgKRebUIS56w1yx5jlBIYbcikTnZH+E2sizM/EAjqis4vYbiZcxRyyPHFwqgm0xqaoxDvYP/
gXVJQsRPR7OjsiQ7tyLHTcvl500zTM2El63S4RTjI3oWG8HGwTGKAZuHSkaA9PTPpnP2vBVNVsuO
li4zN7Lc4PKObCEWFc5aZy2Ho/eTaLHA7wRZ7H2luDa5NckKb4ygb2iAGK9U8U0VWNM5elfdaBB1
XbvEBTaE+p9JG61H9NR+vcw1PYNrMbyncXPINAzHZVFWmovW6X4oaJbpXAuudj9lBFHi2ItQ0VzF
wkzdM32c0COCZUbqe60JGvLTGW28Z/x7Q3pnQGqkRSIRikq99Wt6u/0n9Uw03UqCz5J8T9iu/we1
uB98igXKYnHFRi/eouApnoGBK2j6b1RWl8hRDm9Ds8LXDWMl4uCeSNR3538Jqh13+QTp2bFrl4hQ
mmWvXxN2oOakLKc0IEE99ai2+6rS36lkKM4eWBhYdiwPR6mq53PuuJs+rxT+T/TKKNxDHSLxzS7m
qXGltNK8poWrvNuyNn9moUjRl4nZWwWnIMxShq3+Ea/CZItAkyTwgobzhYyQO09SL++EAqUmIvNM
evsFK/Kr2K14icYWkUJDM4/whcOWmGsyzSugrEjktvhKM3nS6bcQIM1d1fmSSYezWHkJOMVPVxtB
9TBWXydxdWZ+dwxJzbFXNft1dtA0o0Ewj1nRmPe+EOGOrhMDJz4ifyds9YG9ki+rbhN6afOIRA91
eri8d5+c47/nX14XblJW1STh0wVFDQ84uXOOZSSLS8zGZbIn5TUyox1OmkW67gnH/EInbC55zeq6
dLHXK5fCYakMvhwGrWEnUTQfpxGzYII+BSkZolHYs1GZbG5cbjrmJpgY792SuaC9bv0c5TzJ4YJk
kTRX7+UPUkIFvoY08gDS7QIkO4V2ezlShus6n0ZgGZw/HtegDLr3/wTf4uhs2A2igHHl2DSWV2ek
12mxQ6T6iMxSazaQPBp+g5VT/5mgt0824b1IK7L7Hano7Yhpuf30Pz41wb0oklRuQrD7WMkKITI9
pyiU/ir+4QYIWOt+suI4uV7hKChW0KTHXRAuAFjgEqljYr4CahIxnmJz0HryFFLsWG4LxAm78VHU
Jgmv1mJ2ZW+vWHiVti618+XaYRcsmdSCLDgCow1mo6qe/ieayjxPJ7YVU1fSkshPc75bQlQYqW/s
wju1gOaO3yfpDhcJ1mO+9baD9JJEjM6m4wZy5oTKTfCN6iepTNq5dkvfYxPaZptLusDNyqdzwShV
dm4sGHwNiyeIUlZ0CDOy2bVwtarh+KJ139wZ82U+ujJOaQEa8OeZ0U8ZrCmWHL2fcN20HNWdrViP
DRvJL9PaaEN/EKavFUWl29sA6OiWUSfv98e1tsLRXOp8EIiSHoTx/kNgzm1kjV0YCaBdOQvbcz0b
KTne0QMQiUFX3eKvasaAyRyWGTc5C4jU7rDkjksSyvwPgZiDnA903+AfqAxkxbMsvAoILlKSWo+Z
1yVXPPeYpOoA62bX6m3a6wEvJqO8vNLmKi0nuZHHTpTmVhjj11+E4gu/BsmOF56z7zuhR/sR1nqG
XRRm6Pz6V9SQfh81v/49rv1BUK7nqs+o5WEBxsIwmaHiU7Ak631HxYkTn0u9FRmYzwobH65tLo6Q
0Gu0fheLq7Mvxt/UUz0vBt8oAVu09W25VG9PWdIKTU8o7ZXZNRiKYOJ2NBrKiF8XQAZRC3fwbFc2
ecnexky+gY6H8OIWPzwea6RMusgLbOf3X6MKt47pbTPr7RofvygVFibafvDd6UCH6gPMlVxfQFnX
A0UX4TGV9RX66BNffexQV7qlv3miLPtatvBonPKT4ZYKCeSs9i4jskkvrTW74Q8xW+e77GKTAvwN
eBkRnvecEcBFy1tfoY0YGCknQL++EYB2HSFYaWWgf+7UwvfA3NCfZtVUQcGqk1vlKk7k8savluVD
XoQgtGF/pckxlU4GN07HD6U5wuogD6BqDVxlQo6prfgjIt/JcaCjOeQnSPGtnY8Ce+6D/5kUXYTC
HDkmP/AMEcDCMzhsGmFqLD0VA5BAHGupUhI68C1pGOKD/WBWS2kLPz5ek+FxpKr8TswBAq7vkzAA
7S139lze2HG4YJ5xV68m/VBIxtlDqerh4OHSlzVfNO8ZcLe2F8ZI01fP7Mmy61WZztULJCNCZJce
tNqFBClg52n9DxqG4DKwCZ2ZO2G3GfEGj2PakJkp1w+78c/RESjZYQY3KVtfLMnbmpjxP1aYnz4Z
G2LipjOCn0N+PbSWRphk0m/2vuT41n9onBuAZUFekYrzLoHfqzhb+jwYzzpVyC4OGG3EIZnMNOfN
hMfV8oNLpLBYURYw8rDCzLGrJ8uudKMhZMkaOwp0L+vFKu8byicXCzhS4iXObmb3on3sH/wyDeB6
7NfKO0iuXvEx+jfzRpZq/JjtXOpuoLbBzX22twpcBNkrtNNWETYH8dPhdalgq85C6+zmNL7ceSlW
ZqWRgeR/AxnaTMWpawTaposWvJyaccIqBzlVjrbCD2HdsYkrC7Usd5XEDaoRy1jPYbUfvbKL9QyU
VZSzXkAPiMzUqQdwFoJ4kNPAUC/mvzRhYXgk1OuYR/rcicFSG7CVUFY3dyQu/A57SVwdHE0oS4vz
t4l9ulRwuqiSAD9n9zqr1smo2Ts04t7urCBjDM2EmUxfhGXRcYbSwys3N/xEohciUAvqGDQ8hnfM
DQBNwNfoQqeMGU3mgfNXCW6vfo1voPx0W8D44KQ1HK/6/2j7+zY7DOylwrhuogxMTJpBp2MqBR64
oI4h5UIOuXSHKNM1TnUXEgq682ixxys2juB072q4UIvJDrhBl6SleX+dvLy1OC3+uMT++GhgthbW
CTbznyj+5gm1luN7nH3NwInxxMYwGROnrQuvHYQMePM79BhFFvXDfQmqwIrlSnvDBnXDjAD0HmAI
OTdir7pQVQLLNcwItMyQOJSqqRnM+KAKQL/zfYDKJcMeIDlWMqozPlvvLtHJ9xBsjV1Voj7zCTIE
BVcYgYNqzu+0F+JMc2Xf8SS6d8XszjfSAQNDouNSHo0prGAlNcqwOxo13+ph3nnbyNE/SBy22oXN
Sh3Agud4ZF9GwPt5/OwZ0kc8xeWOokE64O7YxTJ6OAP8ieUWaLk/OZbWuEKcfpY8saLeznEUqX33
wRfh6xUGk3YqG/+zLonKLL5hveWxwgF4SqEQmBUv+YVbd1TkEhzQKhM9PiY/oRgDMJlSEAsR4RyD
SEnJZ1C7VvO1dudaJsn87+v5tWRo6DO9uBaBxUr1iVLKaUD1uGx2MhdXDt1dGhXSqXicMnh3yhJf
5KRURDHCxItIWAonGvzj8GpPYcTgkeLzN7G/3Kq6XhEa93364DcX9KBNWq2njhUK1hqxVNgj0YOC
LZOg7G2UWDhYHwMxZh/HXtYikr8oqPKcG+KteBKdqiIDHiJIb54atltH0XIY8xh5YMBGcjiaJUcN
zwLFtmvgq7VaWQKsvyVaTBBF4xMwS/ivME48DPewX1PBsuUiCtzlI7mmnxskxpqHQLv9uxIEHeDG
92aMwv1B3hEVQQkGq52YvQ8lrNmcyvk6+O/DgfDUQHha9BYPvjeuEGKsziYYVY75gAItS3Kcsr0r
Y4c4U35Xgdw0FkhCmqa8j95YIRJc6UZA0E6MPwCOlsYzh63voZIfpWrLR3xBx8B7PKDmEbjSkf+E
6FMdu3AsXVPk81EHJSk2ltCkgINPudTWrUXbNHcC/xhbyGfimnvjhhM8tUBby/z78RGX5GL6At0W
LnkTJrSf4EOyRbupRyo8I20xeRfgHgrlReh+LY+yt6MaEFBVv+a+v93z0JN1bSdilRBYhH5L6i9B
T32FTtiPBg+dN2cZZeEZFu8URDXdpV2n+0Lo8L2INlIOv4Q/Amxp51Um/5cZoPBkf9C+43xqEiYx
+99Oo2vuVM4cAoBXCy+n8T3hq2RY865Tc43Dnz5dUg2Obu3h/1M1fXDT7f5XvZl2htSd4Et8zKGC
timDOUE8ewUIOd2unv48RuwDI42GvDaxY768Fk4G6VEfo2LxQ55p2qmxN/5V0H4CqrUIJ4nSozG+
T2Lp974pYCXJDY3WWLizqwMZ7d6BXQi2mOPbKnL/vnLehMGjxKfeapqoGLez03XCvl+4yo8dkouW
yIxgToupv8FT/ZL0e5U5kjMWKhv+B30/PTDh9QWClwXeFFyPm6QY2Pb+fFHh4joiPEx/DysN4lAF
0I55H8pzMWU1gdGnVk9K7F1OtvsUywAzmzjlA0mosjRmCAcsRuTy3eqdRUpDoZYAmux3pXBHwAmR
q4lqTnslByAgefABTud6sFwlhM9obgRc5bvrvpPU/c0F8RI1LINsieKbUpTwGJyr08+V2kPk5lXr
vYBugVrIJUdC+9sN2F1fTvU5t+ZimljD2p8hswZoEUn/m2QxMem0KdSwtfW8DtJCKVRsqtlyj6EE
eNOq4utXUoHjR31+sr6EN91+ilefWfodjfUovhkYwZomQufpI5VE1TkFEEIlwayzRdcerc/IQYHh
fJNUKW5JXzAsJkO3vM6jLxThV6UFct/MI7oPWyR+ntS4dONIvyTi05CeNDX9wHvM5fAYY057Y/GR
oPVxsyh2Zozd2WALIOk7CdbYBZsyk+Cr9X/wP0uXIHYWvJA7fVli+56aKjXhMvbo9uq2KCwNq8Or
isLY+ZIjfOG7ANi80RZYaw56jHWwbvRmw9KHp75Oy2cy0kWm6mwSXnZVuX2dXQulpiixa82Kehpl
GE6NeRg063RBZboLCS+NKZI3tPxS9xXaX8WG4ILy4DskWJKkhu3rlF7/VlI8Yy6uCBLvsB9kn63Q
4xPkOJrG+zRFdBQDFj0BeoXsJ3LLp0+qRnFDp913rney3QRazPFOMff2mybng5V4TsaX1XdroN3J
5i4u/eg7FCeFWTtXJMW5Tsx7Tru9WW4Q9XiM+ZEaSe0CLDRmA87w2nezZVu1wsgVfSS7e08cf5lY
kHKr/PDr2kwZS1KzwzBPXUezrXOnDaNx+JDKQUPgoQ8K7zhnCswd0LqClsGyB1ex9hldfvMuWnOf
LxcqnHgQHrEa3R15itAYoMZZPer/MymaDv5k3UxX2n2/ZFlLJynAU62oZX//xFlPR7Ts5oxOy5Rq
hLVeVZ10+NpJveMumdz6LSDX9/5kiAqvEwurlubogr/2JwNEXLH+tzUH5LBXfHTvxsmyhQXhTkzd
ZR4sC7n1sTRQ7N0GkI/IKrXLUgxOcw/gUSoBhWjZDxmfU7VJB9yqXsKlPYOPUmRF4Va//34qfuIX
TfCpRsF/eb94g+jj4INbeJrh3sPfPtjqM3nwQkK+52GljJZM/IObNIx6p3YAFiAxuS3KejEO2eUh
ttpctgHGFS8mICD+SgdP3rale3JFa2oqQi8KMhQlltGKDhfnA/rPBYZ/cwtUvO+0uszSFyi8oi+y
LT+ZAvMr33rqXw8tvCLG6KEvcmSfoOQxeCL4BHH6vjRNfAW8SlnrOhIFhUeSx5B8bbgrQpbGV8mA
zl5ScGOQKC2pIXJ1tH2B8W2fEBy4iigqsssRSiflCJeqy9I2Q6O1PNP0Pkw+IR3+MJ+ODLJV9iqo
TDSvyV7okO9hTlnjycTMSbqAm8kv4fa86yD/jb2PEATTPj9n3+qeMuBUaYwMj7esx5CFR9jRa/B1
w75ridrbBOBz336z9v9MaSfZVsKriq3SfLCJ0EYHOJHCeZWdVCfJMtCIK469u2OcBkHWV0i4124Z
7k0MRnVBl+woFTWfML2wsaOaZCfOTBo6NKCF3FV27jdPGBRX3K8awcVRJcULlDaHjq5b+RsOiLBS
U9p5gEGSgmqNR8ummNCiHsYSxQ0puDMScEZKk5uoeQAhm4mqUzWdkaFF7G4NIo2/ZGscDbAqx8et
0J54tXpsfg1qjUyovArNjJGiCOtm2k5lzXKqmkUKPx8AgMhJcscbIWa+pL2UjpYYtB7WvZernGgs
sz04tzcdxHclHU03x3hhw38dPKu2N3+OtentsM42NN5GprlowS8cIR8DBQswFD9HvZlLktieEd2d
RczGHzc8EvF0IUZS0eleCjm5Fqur5vULthKD+UrJm3ADyMCU7X77wYvZrqHKyvqF/f1oZZi4p92M
EmLXXlWVdxT02Pcf+Tg6AQbR4fRmEV7ZPinC9V9Dy1Qt9WS3do1tPvO5gdeGOLBl51vZg0sS+JHs
vJvxQRGvIXMcFDggKqMsYZ+hitLNv2maoY+QK8z+Yf6OAfK3FaX+L0oFnAEHkQqF9P/U/3foCsZV
pBvF/5FEDPIgXNvtcl13ZTT/xvQ956IEryHGuHWuF0t/MTNiQAo8z4kAAEA1LZ9K1pOWN4MYCuXt
i3zV1NW86/ve+GsrlBVJ105y85yaRhzT5R8vIxK+az33ifhk4oz1Ei7lOOTDhJhFiw5g3EDZlHnj
p4WqVkJ6Jum/o8cOkhCmC7dm7wd61S5PCOLos7vqsg2cmAlKbrfuCZJCVmPrQjvOnyeEbnphJkK2
Sjs1C+6BezaOtWJSukl/LTrUoUlRw92VCI2clQwXDS3dLiS6QI3VqXdaGwmxQS8+hgpBVGGyAr+q
bAhUUad4CFYkZ6u3JH4ui6dlrbUvFVud7nttQn75OtuszxlGio634ADS8Jy+xdbO8EpdswnqDUXo
CJtPIo5b9nSh0mYsNs8fCJlMKwS+Cueg9gK8w3PPPmpGLMj9cghG+4xKs5uPWM7PoCwnI/erdiqb
rv2w/b/B/6/9H/qqQ7QO/UjczzlBWxsBo3vLR9GUrvywusWPjG1/T0sFCKIGs540DEMsHuPa4lA5
fZoKTSqAjoPIOy7mLe7abSwH3V5A1K+gqsKqFoaTX7g/wc1WU2yILJKUii6JxI6bplX2uuFxlr7/
j8cBA4jM4PQjIhuKIhNR6ZSiPSkyiMmnnloESoq7YpOn3oASgnlKuDLodUBwy7JIbx6YuvLI2bXR
QAzDDMxd1n4ZWUF2JZmQG6A8iP6f0yhQnUlfmmj0tug3G+nm4PcS7t+3xRQeyI8sl7JXImSrYHw1
98LttBBbwLR4BrRDse0wZz7YGA0lRSP6AzxdFv6VO6u4geo/01sRfFAXJfjhcSYQQjC7IESay7Fv
hMFVAUyLHsqUROUrHO5uqonelzNf+zspXWwdb1JjOVLfx4j/hIuzD7wX+Grrr0TNF3q9MG9Z9XwB
OD6QA+bGW+4Czkyv7HIbyWIzElE4/QniVH4wfXBEVZwjrNwqqPGevyZ+pm0858ueQylAbqZvVFIO
CwSUV7/E5A+j2jqBK5FHQmvW/OTU6PDOGs0T77Q0vkpa4tZkdNnfvznfPvndHPegL6399+aiy9iQ
9QSiK83ZGMi8KfAvLKP1IQgsy7uE5q8jaV2VaMG8TsauipxHMit4xX5KSv7TN2eZWMULx19MByaa
gnnhldJiKF1ZIx1BNealKJupfumwDskMvtlD558mDI3CKUIrDXgKA+aZ7JIub9OS2OP1p4SLr8wd
u9IcOGx0AhuYFjzvMJb/G76dfNouDvH+bFnTyp148YIqaX8q5ta1FwLpe9LnPv/uJFmTVR8M75w9
dWcDjwPvHbA8jbZ2LQji9QTNDv6heJACuqquNwRsyDAHAkXeuuttP09X9W8Ux/bgBmRjtvTdUXQC
80M7sjLc6EqUf0Bq5AY5ii9/6WeMbrk4cBf308AfAoAn/USlBylwndI/Ta5otlJJ1C34ljc7K23o
8cXSoDVbBwFBiaVqVh0faL2/UBNEl1KJxIH7dz5wMIsxKxzxGmoI2tkweEmNbdboEzZp4mFzWgmA
Va4WFEvagGjpjgraMBy4B4XKFjbpuuZ7PKgW2AnFzDPlQnG2fHktxGfhBNR7Hx0Ej7b0dZiYfqib
5NoymGoqsMI6eNTwcj6tBCxk3/XuUyV6UXHmzXjIYST6uuV0khm78dP5qF0n3xZ7djbJkqq2CRnj
Ofmr56VV5cK2y1bYa0quNYFZUBe6v3BeNgyS2iiPOtHOco1aXDHevJ03Z/1VIwAEWm8q2n5Cdo9L
GCWXL9LgPtFXbgwXDdNCj9XW6uJ8QG9yCDZZpcrVVsKDbOouBx4Rmgu+JodCJel2xawQmbUi5DlD
QT2MaoBEXgSbv4li1JQRyHm6HnOzbLhQtEi4/49Ss3yORkEowLvg3erAngFNKVCftYeIF3xjEIEX
cwfzn6MVBtQr4LLcOoDhZZFH2y58pxOW0d2nNiM4upHvIxHBwVTKO/Uu9m2F58fEpqq3J7C99cMM
4UWt0r5TX0MqbrpBK5kE3p/n7wwsuhhjPVIK7OvGQHYp1d0F6LyNURN4iRcKht0iRcf6T/9UOngi
1Tp+cRjDTnKuR/1g4HTqgt7dHAnIdrpu2zErzuRgWvOvrbGHqg9S9LDmvVnvrryd6KFgKPxt2bb4
CpSm1hYgLf9d/gcR1xOAv7cE1a2UxXCd0gYUUNWaHgCLpGEaEM5rDktYl/CJoYdrwdekUQdGwUaS
pc7V2HqvHhh8tD7PEOb91qMwzRkwA7zfOdQCukYdgA3/HQnnbIOfvORunfZdwTeIrVIwZTHb6xAZ
zdXN2anCeluGLP5X1fg9lNn6XM2uS8B+yBY6RiZEtDEfWin0VX3cZGt6y4YzV1GACWloJ247gPat
j3jsxJJ5Ua+F1r+CBGAIDO6jEzhVJZOZ0McxuHZ6QdDvwzG6ryegOpVov6U5a9GUuJz8dzf32urH
TiO4JA7ZHKjwsRt4mwUjcOCLJl57A3MbTYsYpn57cWDMq/93tqb7+vmhis7ix5EXUuuGUoZimVkJ
42oNhEHfAugP0WJPQVeB/dAtSaKankG5SJ9IhC3gxHikyIwGe3q5ghaO5vO7B81ANbBifg7Eres4
Is1R/Uja2BEacXbwpqZATl4R+xTFb5aP2R4kQaTyFfRuPFkWijcXxxVkXAtrFthrVU63b7zPD9Be
6lBJogCuR+BaQBiNczIm4haKTz5uXd1eXGbBo9HyMvpIJibVci3CZDpw0UBl4TZ6fV8od0p7+i4a
jyOWQnx+bEmc1RT8eQcgaYU34wdCfL6gEWXQ7Jy9KXhOOP8+fsOqKxqcNNOPkit7fNv9zJhOzK2K
rroaP+ArA0/P063VWXMS6Uc4+CG3U73bgRbvZ4+lDMI9Wd3gjOxhGy72vNCLTNle5/xK688PGj7B
yqhi+OZ5s7TCcmu0Ll7851f1CzdmwE23N/yfxVSynMouGwMJXJyzm1AB0uGTUFFgOFBloc6I8zKc
JYr2Ucnbwj7bitZ0n4DsZPGBqfIGKHpQMe8zl63DPKrS6C/p7na6bAmpBDfrcouGsN13bRCQ3L8h
0PeClKsESyylIjDJicWtZ8ByDIiX3LiE3eFGe+j9xq0L+6vqKcYzKIA/C3Epz0t8HxtpTcRVWLTG
xKZiOapRN3eFjc9Y60pH49VFlQ2O5ymKft2r+vT50vWbSr45ZINXo/SjPZL7JWPIAgOX9B9x0NYi
6uaSsZRAQOEy3SoQnCMwFq0QOS43n4sKGpr3pqQRrgHu2JugVUnDmlR1jaqbtIuvYvAVmSw6sQZY
v0LyqRTD31G/sWdEwo//xm0DRR+WnytUjyjt5dBi5AvaNI7d+Mwx6QuGU6GUQ7Th5prdSvaDr/MM
nc+IxD3zubJ9pnvVxz/BoRfoJNL9DVfSDbfQYgPeFYGBK3T+ytdo6Qk51isOhUFeTQZj/nHYU8Nw
UHafY7K8ZuyqLEqRWAfPdbIBQuK77Y4u3aGCgJ9ohrEbiMKbGryhPHRnB4OXcfmS7uTl6mTKFnbz
6XMmQ0Jq5xlYjrQSaj1jmb34O2czDUVTGic2FfjuKCwCNopcCJMX0XSOagBuEYLGx8prEGwSryUa
LAW8yiaBHQ8YGznrOfpYxkgNaPT2IZGASLt4Y/5by11aPdoMkZY4LJf/qVsENmKziMVe4GX/7zV7
zeJplID3Dow8C8tGOZ2W5h39/onfwNyEQw56WQKSJRzIa6fnSoouUsaVTizilh8UiuYTjyt7ci1s
tTVsnYC+O04B9vMOaWlG1Rpm79z32qsjp6fvkv0PLEczdWCBuEztNwy+Y+A5DvBx/21CRUfi6I+x
yCQyyIkAJ0b52Y9kYOZu1dip2eX0k+6z3gyJOHAwM9O8VSssvYF0U+zZbj9mKM89GKW4VVdAEVBz
TL4IdHB3UUU8fmFy/HwaTmVYHwzIy8fGKwR2hiZ4yTjWswcC3nyGwXL0opu9fOaV1759Wy2zcLUY
91ZkkQQb1BFgrrzT01SJcWISAQ6ezrc5KXzD7MduLcoQa15QUAIkVhb2yEkW9WRdeFTAtS2td9oG
OV4/NwgvemDxuH11mDNTJyj9jMwyT1QDbNeFW44fMr7rBJIIoTbGC2dS7r9BKnyxUuuCvxrpaoVP
3M0xf/+hy6MpDwxRFumC8/zuSQkxDFxZKMXdmAoixxhd0V1otxGnPqkS+9tw1YnyX5F36Wo0ekfD
yuG85t0BlbdhdqH9VvI+oc5D5X1C0f75TTEsQRhfFdNcIFPrt21HHHsIeZo2lVctjXRyYOrTxJGf
c4QR6lONIDuEUv/jOOL4KqnzDetYHoaU7CIH4gsDA8U/+U8CTSUIHU6Odu/6/VqLGpRnoHeCxDSt
QJaiC0UuUrQyF2T7+HElphu6/09tY8V8Ts7Kd4I5SYptj1tb4ov4q8oOAJIQz29GMahBoBVBW7NQ
H7g2gNNzAcmAtrTeIWOQZ5HFkMcsETagantaqHzfSWoQqezrIl03FzoEFMi2eeovUWMFDT6EMgjo
S7kYkiI1RuObmfjd2/bKThyeshqgKOtUI4KPUNWqiNhOrQZE3YsXrWj8VFhA8ZBoVUkNaOuEq1cr
tKnoDKg3+0TDbhUZQIINoMknmG4vXwSkFxIP0PtzQ7EgVwezNc7NDRSNR7gSfQkBe4EgQivmPlQX
fLg1cz1pvtR/waW2ulPx4S4BMHx+jTE8+jQiQiI0llJReKdFd06XJlECV7GNfwNS7i4wBSn2aRul
XwVvTc56NnXlRQkm9BM3VhzHoCk0o1WxilD0QmqxQchPxE2fJMiKvepUyI5v7qxMtGIiZBXXRt52
Y4MiAUZh0wSYm5EMSF9BjJ3SmnwgdH6NCaFYZHvFov4hT8yYzqpsOe2ihwx4aoKP8zi4mQO8S47s
negvJmJILXXYzYuOlQActjG+3vuK354ax+umVerpKLbOCyeq/zXknPQroh4nAIgQG+cnLCMzCuT+
TD7acdm5SRMjAq2J42tULVM++SG8vTgdAQF4/qN5qwZvS91g5LQdTqt8BAIew2sAPShgUagiLaJ2
0r4wgInEDjY/ZBPtrqmI+mijBWxtObp7oA6vfPwMb4ZUrWy7tgYWJ1cOd6eyui7t4z0mvPKFwnhs
Pcq5MWH2aDFUkQv8stSaKphcCFzO1OD4Vf968Du+cabbXn3NrxbcV1+MjIXe97uMmm6JE0p165Py
Bpxz8h/8DVwyoJ8Z0OI0S6024qlEYEzRaPUYJTetyNGCf8tYe7xUbOTJ+62m9cG80NqlpC7Rini0
uGVkgy2MqQconeU2A7X2xNWhEMINm0vUBF2Nil2qO8e3IoO7NJwShHO+gVbOovCOoOMaTQxcFrM3
5b+0JfMUALma5rUhjWyvNb3evCuNNMgPyn+Q716Lzg9gfet2XzA5VEK3jPom+maIIjdOcYOLrfeO
NuIfwtG1Wunjo5T1x1z4PEWCz9Bn3qq+uSQ5P/YemVSb2B2dQe+ENPP/JqoD1MD9ALh7+hzCA8WL
Xm+Zj/gam8yeu8PL7txovA6UkKbnWJuAj01BQ8kNBt1HpQ7HEtVPMMpfEGv2cxJRPAPgLdZFw6on
cpMW4FIDtGUgqxvZYhKLYWQ1ic7MPXOTQ2FxN0IVmJizpASj4H7AuGxkhBPg+iRMLHZcQErJrXU5
5R9uEl2wntGAk1bJhyEf1PwX4L1e8EowS4Wj+FfD8U0K3YyVSK4TDJFQe1x7TKTLKD8tWAFqFn+t
oocQmbldKRJvxbLCcf5b35h0zySD7DlscEAq8Vvx6ReUz2wSAFkC6qC2SC1Uh2CT/F1HSAPFmBwJ
zKFEmtrK4bkRkb/a5dytwoLHype6ck2EgwdA1TSC9P1LWoY8KPjFbBhG4F87Nh6Oi2HODBTDBCFD
q2oRUHdNZEOmIOKNihIlEG1gFC13mKsa/BsbyWpcqW1VL4772jyYLVpiYolcJfFNCwL+b4/55ZSX
X3ZgSbaQvAi44LtC4M1qL1MHuZLFY50OnKn6VN2QhCWvWAI8bnDFan1wDvh7GvuAIJPqpOlRvA5S
IrySW3onLwyxsWOq3RsEW0v47lVOMEM4UZQHEH+l701/AWglkJ/Tz+1qdUkwYwxNXFVWpddz29XM
kRG/0H0aGl/hdu48tV138nWw8WWdh+FLuu5+iiR0gvCXabHCexF8CCotdrQvXoG8gUQm8QMmbGGz
oW6bbT3HCvwc6+3ndYrHD3bUMukz1x6M4+H7LpB1/lpaqr0ldzaJLDkc+I4q+qL91OjMAXSvLjLg
b6YwtGHiEhFyp6ZZlMpBqwr6E1i0LTY7ZujG+drz20UKVG9JBqXsDoUPidt9B094mYHXUIHJYzAt
RlLUJJCGz6xFxbY5NUCP/Iai6O9VdebU/5ryhe5qDTxYSRJDlZSIw9z0jtZ8brENlVFcqDFiB3la
OTCXFXqoYxuhf5adNpE+QorZnwP5vfRIbazmC5AjUCnyIMXqrV9b15gcfy9tXSBdMHrSfuzmTjvw
D4WhOnQ2ZDBc0seU72OHnE/yAG24cgkECnaUn8n8q1w21rD/pHGNTaObkDJ4NXlRnaHWIaS1mRQs
+iM6D5R/QJLvYxrNMn0v4Ml1neuig/hb8obAlYj7s3+TnNI9M9LpTFlN9dga6KtbMl4fxRAWL+bA
vYCh8DrfiG9ZekIyOjfoQArgf910nRZW6gAgr96plKpIWBrk9YO6msvCXiaEgpQQ7T7MhLomMVjD
3K7vIqvr/0scDqg+EL/WP4Td36BO6SiUwlt9+Z6NASBQw+z9yRqWFHrauVQrZLBJ/WISh//P60b/
8vteKbCEF/6cFZ/Tr62N1ZYhkHbi1mWRv18W01CAsVsTV05UXhThtMel3VZ4fhO5OJ7eUP+8q5My
R1rtmfcfHEGiq2qy08gv64XcAcQqeT7ALOuJLMHpmA7BVoJeS6QnsyXmr1UiHXSEt6CInU90PCn5
KOy1c6tD/uAO0bFEzWIdR5UoE17FhelXbEY5JJ5PmYGjPjJ4KMKonfXg/TCDbLfT37lgVNhD6VRw
P847wlureDtBHK3ODxKfG5qMm61F4U5BYrzjh7gHRS3DPk84nakuF1wAgaIuRROp+BUDsjdM+Di9
MmvIwbMLJgBZZTkw2Y2f87it+ze3+PsKkpVqByYTeCObYg4+Zj4aQxcl6N/HLG0oKdv3jgWVUW34
FI0UuDyWw4gFelo5VlaTlVW4FwX+CkIoKK2UgynkP2T5FhTn56zZvdDsEdWcQpUv8vXCxXFh16ao
e2k1IMQ+DBZXP/RC59XHPcxnOYFikCXlPpHfuz6yBcnVf88zjmGe/0axIkEnUy4vHj6etKIyKuXR
nQWyM8fv3sC1hCyrbjlcGEAqG1gQVfizBTuAcRI7f9W9gaWy4cC1GAPJktntU0UiW8cemGqskTF7
XguRHcrvqgKzgm92WKTTxSO7WPVSqvyNsD8FrqBHYvzPcFcz0muSvbQKj9I7HGd1d50I2lKZa66O
O6bDAcIPRDrwWeHh9RYxfZAiMk44Ttbu2SMBr8Y5llM5gTnamY566peerAv/nBfmHfPjJ/Ga+31m
JKcJo3ueJf6IZpgILw4zOMruVFVesSKDxolZ0VR3cQTc+hSqmqt3T59CAUULAeV7GT+CHxcQEdYT
aLjj5PbgFM4eKUC3w0Eu7vs28rwifYj7xNG97Os9rpspvWLiAlo9Rq/WUsw2ypBNR6UxwXZ2JKWQ
/ksN36t+Tc4Gj+VaMuvMDlS9hHELtbAEQCw68pdQc+/MrVnBD+/lInGGZd7+wUf+3MStAeukdcVr
uRZ0WnzHJpDaA8i7M4VIRsTiRfGHjlbXinTwbjvgd7HeBSVWX876ftdmkUs7yzsaUI7JJ/q/GPiv
h5MkVMPyRJVWs8K6R1g7WQPmktRq+/Y2AYataT9D/7+z+kWCm2HAD/gh0vBxS3J1W7UnXReN4J2o
K0Km9H5WxWZ/ITVRIfNpoSrzeu81jEI2F/mrRe59MpldH7QvS0pPOyS8EP7ME3mQVGdHjneZbZq8
rT8+OrVzV8hkT1IJagRrYt6GWjb0bOgdWUZ4ogriZmiv4ZqfDPbMkP6f0XwbR6qhLM5PuLpm6pos
mwr/F6HRXvMd9WlnYRyADWc9sKURwgVYrDgTpUCEHnQTbhAId+0UGZ0A0wWhVl+LMzgLJpS9qAoz
KNYCPFJWW8U+33bYD4gu3+hXpbNzidYvT/6OvvcFo5MnccAboq53auG4R0fawFIf9cJ80KLyhlb6
sYToDqYb2NXcdLICmxMuXes1+wGzvQn9XBKBF1j3aWCaRjnVNvVF69/hZSkYoCzf1D/L3+2x+jBm
8RVTbFLj4lFMlC+x+paao7SuFz9eqNVObE4N4oXM8HiiByIufutCo8WvmsHFaIJNCcXM8Yxi9dna
Wz3ILt9b9dEPpeLSRdpY81wXi8Lnn4nm8xq0bFtkvNR+MBXlALVFfrGcCBPm/odPFE1YQncT2uvY
4nWG/wAdiJEAWjIbv0qWrLhAaIO3Y2EXZjn8Fs434TYQcT9udR6DTEY7xF43mIIUGwd0InjqtP2N
Y5VEcqya8f+9ZbqNUf6oWUpPS4diLtCwIcRvIfZEsa6oZhaitishYMzv5fd4R/RCT0dbMqLYvU8i
BO43oLkxvYhVW18vwZbe8A/FyT8GRrm9pPGtVmGNNkjt6OL7bbknTXCjPfykQ1wV6al7Nimva0IA
ZalNqIEEc7bqv6LVhuczClLwjVYVqZHQoEt0mb/xzM2AfV0eJkfFELp2sdb4um0nFb3ETzdF1dhf
umxAlUucswxfDdxeZKAlxLq6e3RctyiJDhZ2UZuLj1UON4roNtO6ft/jEsgalmu3IJBYuN2a7e/3
Cl+UhSeKqYMD+CWbJl5t/nqoB71assgWBa1c2EAubvpBp+cNFQ2TExmdt4MnzmeEk6h3Pe/SvmOF
WYoUVjB86z0bAU36pjJHH/0ZDXboGtOGsSiOVqYETIgQG0Mo0G1ZaMhqOK71cDIS8uiDfNnLxyhP
KYI0c6yR8ZugfwIpYL+JXtuW7Cc/3GmBUeOSiWyGjDiTEHyrBZpiOoG1E0nryOtlSB2HKwd8Rj6b
2VLluPlUkDjYTffZmPcMj9jmpL7/u4T1ZPzthEpCo8CiONtMVLTeaMzk+k8iOGjr612DZSgLr5MN
qnIT+vrgHLyCFoDsiHmxHBPJg4hBlq/6FnMrvoJQoz/Co8ZRWax1LnJ3pK+Q1ZlAY90OgMnbUSj3
/NbgdA81wowON2R7EPSWNR+YVBUGaEl6JroRcL7JJ94pfktrnaL+RrTmtabrQhp3H3lLtzt2SIAx
8TF3hXsYTFiALzPNwEPa5x2rJhX6OKpGV+YG+ysSX0lzuGcVOF5VTt3czw8UUBxTCxSiuSWoGd+z
szBkugHfi8PgCF9EMEQNEb7akchFYSSUV/OQ+haMJbpoevH0AV/ZlWfQf6nbxalr8Vcuk+VyaiLv
DSXgkYODdtixVL+7fgwv+xxu5Ic9mqqt3jgZwlZFfOpHe3OD3EHYUJFesZmqlBz/7XTYUw1Vy3ma
A5ByQT3qrZMp315eMRl+fk7R+SzcI7cfqA1eCIp6rNuJwRWi0g1gx9qu+ebIGTfNeURYhbt28uJn
Pc4TvlZXiF6+FdIyOL+AlIT8Hr1ZFYKlTG00aDzZtVFOCP2CUFvFkfYGrmhSlLSnIxMq2eIowUFd
sxzm75/XaDyGQjSd+7/V66iN26jykZJ4gcjFQwMard1txq6JrDilbZ25IQ3w9B0Rg25zLJ2PGtI+
hUCvzQBf4qEU3kdEGrUXaXhshmMDzcBzxDrI3my/wfgq1B8o0n3zBe++ESjZaagFqfcRi/kRWCtX
wBsO4DFpYHqOqwOsuszzeDWSlsiHra7TZIWUnSy3a7jpK6Kd9KJIueZc61W6Xt8FTOktwzM7X/dL
81tt8DtBRkNODPgZySxjlg03OPp2xjY+MZOk04uQvcqWsui9K/ZrvqAZgolgn5WEEXWWQR+K+O8w
iOHBbYRbr53hx6J2yVO+JVk16F6nCGZGpUtLWlKy+kgJi+soNcdi3hMisyf+I14kY4cTSxDMB05G
PkbEHkaHSgjZgIimyuiG1YVo4eG/koXzgL/XWzwD2i3VcH2dqYdEgxdqUniLVzUqftFgZX4SCoiu
GxBcVfxdTZMBkBG0krgWURYzWvNwZ6ZgHLC6k2gAW4QWIUhC+1v1s8IZ0CgvAHV+8DsMpJze9tFt
VhPHxHWU1t6sbsbV1/wGJirp8K6YkW5FlCqe/6Ha29+W0ohlVlkDNoSTRCLBaVq090LdugpBzQfe
AsJOV0nVeQvpOZ2V3dU+MKFBjuN5deEY39BQpyDPFpY46Ivxn3nNTYNcv50N+7PrqQnBR1BxoDaA
ArkQByZQBRTlDk64VSdZbAfdr/J8MxTdP19Rf343tCo05R0K21U5Uwe7I89+9KFrztA894M062Yv
d0ulT4PtSxGTjRqpT/Kzieb1vZGC+ouRaTgydWWnBImZ7pP79HhMIRbgJropRG5aW+3tFhXf4HBO
18XsYNLLnftfB7Ibff3v/JdwDeI+gLdZ1iH+00J5TowiP7qE3aXig2xEinkhzp6JsZq4iEDjVlmq
L09Hla2Vjd1BUYnvdp04op3zg369CTutoCq4w0uP+iig5HgMRebQ8rXzFKpv0JsJfOLwkf4/cSaJ
Bvp1ksqi2Dl/SpaLndCYjodtaTmsCXO32nrVtCx4Pka/ZEqwUbf4a5NZriIBkmQySNHfgYPstsIQ
42cuSUeWncAxxX5WKegdWbQ0PIuh/qzvoip8h1ZR44HUqFjUsRRXU1F6nDlgZwCPVq5T7taF33xa
RgbffEJlHpD7a8PIpW7xitpVC19fRRjv5ieQjlFLubJZDDH20eW523OeH2vkp4TtzAtUUkQ0LkMK
7wQ83qq8vGp2dz6SaFVHYJJYMgVUyrTjg7k1Kl2amfzN5mPxZRf71kDn1c+HTVLRxz3DVeImLeV9
c1dh18vKNK7YGTzsxrj4pcNV2+AMtZDcnAofwFRXUago/uvCGLHqOHNqbmYVBS77Wly3YZ25u/qT
Vejl2JQKC+sMuqyh0vRRyaYzib5m8ZoVeYL1kBMClxI64VYQCEumSdedhgCb7/Wrw72bWTpf/GqY
rAyWf242RKQm0BKP8Fmz0oOvZ8o6qRqaDJ5IsoXGvmTyNX8qFFay2xDdofcIXVCOCNwgz6Su8GZ4
rmf8xMPw+REsDPMwt4F2wFnOqNZwnXH2m7IG0bMA6cnZsv1L/L7myUCCpGxoh1jM75FWmbvp2t9M
T4HouxH0MgU+XK/G23PwKNSrhQD7Ur6ubbNnPWTpkGZq09PwagVf5CTeHPjXftDRbvS7W0f9O0z8
5m7cgzb7+aK36bCDnyFW+2FHa20elnG+NPXQy3f0Wr1Qq0e9Ho54SatomZfvzeph5WUkt5nJQZZ8
Ybi5bqp2TC2uL0pl3hA7NqMnj5xJgTjphiwQig/gqDGBOxqxuQxCoyhvhwqFcN7e/8MVyZZFlK+/
bW6ndX9TPZd8Nm2BulqKBXYfb8zHOI0OpHKAZfe+PqmhgF0pAwZvZZFVAX7PR3BH7EFxOxwx0xrD
DsGtf5UFD7XBSyJOyVSxeF0istQtVniEbdraEl5LZIUUstBa7taEDWN7mjDKPhmzWGF5vsXgmL3i
yhV6+ypNBC8BGLqsTU3zLRp99Ww4Rc7hQuj2rIayM2ClKQMCcLCAx+fWd5xpMbzdBbyXyOxfRLe5
D0Onv2vx8HsLBcIZSQZ/EJXlvXL7SHIDUP4nWn/EqVdBhTfsZwrmWQV9gxnOxxOKNKv1gPIgb2cL
xkmQEEJFrj4qnn47Drp3CGFUmLwfPXFL/4Pc4+cN/6zIOUbs6v3vY+Ljm6fydtfnA/+bb0xrcGPn
5Obh+qaBTsFMktPeShaVX3v0NggcuY85YPjP4HeHrXn/OXOE2GToqULbjlkKeWciHEZBCcJKbzrU
UhF5WI1BUBAnsGTI+C1iW/TFXvXeBZ+Ue3a9MD+CC3DDauj+iFOlpMIgfxzbsl87q1zx8fBNLeCw
HA2RmHLq2iIyVLDLH1p4fiVSZ5UqehPziV55Q1G1R4dIJU2YwJvfrH/wB/CEL13sPe61qNaBVF+S
ORQozMNZLBofNdf3QSi/lWAsPmTxXfv4cifKW6OcEbdd5SI1i5YiWTKiJdQhAlmURFds2093FoJ/
eIaNULOqnPld2D6HmGCRShoyEfVZhdmBfA0+w+g/vKHQwCKVXFqi3DBIhK0f9lRTk1jbP4dl/2Bd
28s3J8oWm1ZaG/0OkfrG1UrzJbhlAiyjgYvNOJQeD8aq1USaCEUBoffAu/XucFRulVaGfpnOuLvZ
44+B/H4Ku7A/mHH7usvbpTpa/2vf2B4HlyxEuR/heFRTpsGkNkZ+kvJdIBJw58cOKsHIuRiGuHDO
ZTUrjS2yFCYlGTNZcLOIzybyBxHETt/Det9qdF4jrWiGScJsfXM3HOSzeJG2MiN+JwsSr4VFiwJX
rY8w0QPBeuRfjZP3qMCXfHY+R+uVOPuSMMOun+z/l1dE3VNX/vPJb6KrNKG8EWvSeYLpxhQf1dD0
5tbkaRCGNJQrfYzmpTHhrVjdTAzSubepFVPfBj77PijH1AG6pKrnOmEMRvTseHYYpDi4+Z0IOysi
bU1jTLZcURBjFCypY+R5iuZ9lov1sFic6Het5nbnMilKQS3gdZFONlGFRWKs82UQPLEqeMZ4gWWK
kOkMbL/vQ8hIez7I7djSZRNpFOyfwxMlQARGV0qTm21Sf5BLPY0+1WIZSfI9+sw5peZFssQIeeMl
+odzsQMzkLb7auqWssIHXo6MkiwGRmrfVF0bp2HaofHISj8V2OKyGZn5Kt+wWrkneY5nQ3B+7w1l
MfBDeZhIljhAMDSbKG8rHCXcyX8loy6C7YyFqmp7P+MUNlvO7VoV/G1KteXxKBXdeEeHyMP9Sjaz
BOGpa2/nGnV8aT3Oxl0czrT1Irj7m8ABNoUXKjqwbAcZ7HdDjgV+UDX8q5biCTh6IxdL59S78ZdT
j2P7H5nni0n45zoFzwzKF4JCbS4VPsuaVpfFOHh0BWRmCc0L2kv00IiEgDuwbZPTN54UGoitmXgC
f+ChrfQr5AKpl1tX18QJpEV2QzZKsGcG9FZrHnDzaFx2zOV/rurFv4Jq9ic2ISKNbCrXud7YiZI5
tnOxMN+RXt5S0NxGaMyhzVftVsu8QRbOWyTDmmMseieTNmvB/huwyoUPJgqWDky+NmpsuXiYK/mZ
Bpi0cFKf6yV9UH/o8jtt1cdFhWdJIWqklMR5g0gqdByBjVQo4DJf4liwoMP8dkz1+CofUQLUcifs
CRdLyAGKP4ZUrRS1pnuc9v2OM+9CyGrVlEgI967g8+4ORoizZBW3BP0gTWlnh2qG37ROD5MGFq4i
foOhfmLdNaISG3rxygXKGRRT12O/aUHAFbPF52irX5RY4GiLaGG92/AtofC6sVIHkTFtqBk9vsM+
qF6nndh5iE55xAX+tSgYPf1ItbD6v67cZ6KFggsHxOoYtZPwOKhvkxh6HVZRcV5ieDB8LVFS1Z0E
rfDUub/RTEFtbAOjXfKWRggLAaEmk5250ZxFWNaMG70QSOAY15T7650LaogxL9z42JA3feg25L87
OvZ4rZFcCq/9Trhk5W8Pf+qWci9kiVabNAx44ECsXcXULpCT6OGdO4rs/7MeqHcOlGO/x7pPlXlr
81CqNSgnkLgkEPo/jYwpeWPBAmiJHEfjuSEMTHD/Y9ToUSvR7GF643Fku14Mfh6WtVwSbh06vD79
nIT6N03gvOp3pmdhfSfw8k68XQm4r2a7CXXbFGm1N0Sx3OEHCl25WDJz3aYGa1JBiMhfetY6nn8I
d6igu4kG2KB5Ir11Hue+IoRK4MEJ9ONZ+d8MdD5GGSHT5215zyH8aQ/deBKKMfzja8V7MHEDvSep
oPIYJ4BY4lLq2RtzGWxx7PJoEEFnKyf/WtMSx18n/REyTtTNa9Y+Ws4dCcRlmWtZJR5uuK/h1Az7
Lk05USEQ/jSw5Bz3S0URkNFX+AxLCJxcHnHRRyJ9xW8h7B8DNKeohUDxFZdKXLMIaahqsdn4SSZ2
dN3IIdJnYIe9F/EvuI/1dFCPhEU06f5Ag7mEQPns8tvPz/35twEW39XiQsnPN8yeH8lvYLg0gNrx
FRPOZRbikFBK2Jv35SbS9i0O6rJvo6Bso854jpowNYyjU8ewK1pTk4CPxFX7CyBE3L0k9gTGAsVV
Y+kUR6BbWg2z69BAFE0lZ5gXlUGf8uSihSaDZpv3ks5QxTynEo0701moZVpIdXFihOnBT2JIv3LT
B0l/L21tG4Rd4GXA5XdgUHtyl+Y9mOzh5TLLVGHSSumVGRhsTQgkrzslQ1hcpmi7AxldASXEZ3BF
9TFqvaYqZsQWjFwceE+Yx7qQE1Z6gJqihZCoKr/LIqLjlp63qsH491aYk4/uKT4vMegGkzgh5PTa
NTIMKY0cyxfkvdeI55sXIhe4wNzQLFqLdf3bfn1jrxiflco6ZAvx4nw85YQli3cgxfzREYAaWekz
/C7quhKOzWZ0uSBdr3wSUO5QsxAYDC3BHmnxuJgSc22LaNqZSTDbafSTIWFg77plk92CVOpAzFWn
Fb1oJtGRVs1dVfLCcMPwBKCT0xHH8be/wAkUipPTliPJAsv7ZOJoKM2MB2hXUu3e3yjATuyrbgvp
P0f+x3m7caS3JyyFKaDImLOCXuhBOQ7b20oqTgkXuE0u4fBhTtu+VCdQ4fm2YlPQPj1LnI4yllig
z2h4RN2+ReKNYzdoEbeFimPHGE+dyKmZ3nVtxhjAbkPz3ToMgp6Y3WV+PPW7AQfUbbYmjh/TZ+3P
zsCp6F7b3SIfgNb7GJGtwbP7Py5qBeyJm8llkw31WQKDaOzus1uB65xRd+M1d7JYuH86OTN5Q4V8
UB+8AVtKXtKOVMXWxIbRgT4v3cz6Vvtwu2mvqFyB5ztef4BLrh9EkAPgMEDT9hIuMDIscgPmP0S/
+rCyf0f3xdsI6ljU/ExgW+bnQKBbNyZxBZt7hGZA5tuRQ5Pnfq1/IKUr0KeF0MgW0PnL1YXB0tsZ
tA9U2iXafezmahQSxD9/6k8CsyKzBbxX00B6Htc1ZZXxbW1jcOPeoIjwQP5WVUjoZD1NqZnYAeS4
/wJae9pro41rcxrjih3OoEcimo42DZylNy1VzoA+2SyaAju5tN2AveuXVB3NL+aElJlrE+8lyUuW
fQ8a+2JTeU+iIpxZ8mPXsfD7gU3JMMA8G5F6+6KkzbFyM+1QKkClq1U21gCkVx84NvE1hDuSVITJ
zkyqAmjF9G2q4rc5L3NY0r2Ype0qwIgz6gcKNSLtE/Bqp3mSOxiDOWbxj2cg3tJTfspLuTCFWLH2
Yw0zhI3AioozrWiZYGm8XwJqsw9lxj7FDdGNM2GTyLNQMr17pudvTvnB0yfhmQUk5Jb/iaFb0WdZ
xy5cWin6W2/26fd3sfDgSaTxd+sZCjL+puLwAV+DV0abd46yAED6oPq0AfJVBbJQbyuNA6oWd6IO
g6kDs7OjOJYn17CbmujcKojNdmqLRIBR17jgZTHfnkDQramIuptWqGxwsPTwd1y6p2pxQVrdYdCD
T4hC5csc7V9H+63UMJMiEOcJ1MatHrbqMOH833Jh3bmtq7cfys1ZqI7emii0FvWY4W2kagZdYAjc
A+WmYxMcd/ftZMV8+Dlr8mUTeoM258qdwWfYCZbAsGEqWkAARYuqLmaiWu6iJUbBnml2azWKAsKD
757eG9bwB925gyBd3FdCUvZf8jy5Dfr/JgN9rccYrPaB0bwfb3kTf2HruI+Ax7SCjwQ5vf+8UD7e
84jMQe++aGZAf9P+5oWyxP0WuWeDbeBxgn4Y2SMZAM4dH8wiyY+cKuFch2H0wMWzR0d/O5UqZ83a
FweJPSV85MTyodXkAj8LvMkx3PAbndAj9dgs2JPsugsL0HQE6QWb0Z/nQOlhFIjPAJF/Ys/GjPAB
lNFhPHSkg3/iyeBmVIng73RSZCEezmvvyarLh4xHsBU3RAOSmA6ceeC9+uLk4LyqSIkuG5BzswyI
Nzk9cTCTi1u51+QYVQJuyblpokmMJMMCVvZbUmnh5cE+NrvxoH6JFG1fRqmbRY+eIVyHw1B24Y4H
FenH7h2DZQNOpOvpTEY6EqQOh3225isHww4w0rHiovpbRKelZBfBKMnHe5ARJCkl2j2OZipDkPCN
C9gxQzRXMs44gHN549VZhXK77AJm7hO/WMIwMccideF3jI8rTkDQ0rYomsnpjfgzZCuGm5dUkitZ
U3qYsHOffS1YyZ/tgIC8+lWRLsY/KlaEjBA/tJvAthb8PstWqKy7Irvp5KykaCKweiD9+4BmRf2R
Gbv4tcbG9k3d4Nnn6TXEddzl1UskaYcReyTFPDXFYu1PX+OwKlENP51LAuQXyXdFf8H+6qIttcOB
SmJm0TgScePkV2jGAGzIQCrDgqP+5Vwdsb9dChoDcFvrhRMNdrCIydUvZMd5fwD8kFAH+NuLZ/ce
vsVQfCzQI3xsuZZIJmhEBCoa3bk8+srpYCaTMVewAGvrEouY62ecDm+8LgYciZLSPMAUJ4Y7Ur0w
NE8q3qeteHHbw1e9g4cCaczGvQ0lUTdOBTIpdRXrEdhykCT/7VYJgo82T57ptLW+BjSHFRNsgE1J
ca3+Tx3Fx62joCCD9OXWq0M05UaQTprMsFt4AIyMV1F/MNROAlQsIv4KYSmbvuMg6lY9J7kXTfIE
wpwefwxUB+sHu3c+Hzs7oT5pf1nNsYJQxqnfL7GEmZZxk2YqMfNYv4FUSfalGmd4SAuIPE/Qx0m3
+QmYLqPePYYYqLLQNet5pKleoQmd41W2B+X25Q2+i6+VHeX0NHfWm8JrOTh8daPYrcetudPTQJWu
T8OZhjfrCSabvITC1lJ2cFCg8NTlDBI21kYaunr6AYxqfEVOlzC1KMA8urVuD5lXlvcpP9xkJYAq
H618tDoz3savk6X1baduhtDhVXRXU7DKtKkxRqZsoBC6XdwAcxd5tS6kSqdCPlMAIPnb0PQOrZZS
Vg2dqHheEeGtVG2BiTA0Qfm3HxUVFY6Tg4ewxYXxGhXDrhmT/hwvHFDRfLWaou/tNNIVymtKeH6b
naLR7GQgd23gLXBd6wk+r7NodAn3uC32x2bkUqL4bzjEc+E0AVW2QKJrrfD32YDbP2MgY6Rh91cO
zAZOikqumYj8S/fGgt51cbUL2QnALpZgoAOKnZ5VzjQVMM4KJtY5vEGJwldTP+B6K/k+tnUTr+WN
DH2ZDTbHwZtr1559mWPX6+jSBnnMpzM6IxBY92g231BeBhkKxwoq2JmZo4HOl4Ayv+PmYTKYce1e
yRhjRbeWYlU3vTXAJER9CI/J9+BBycv5PVRRhnKByoVrYwEsKH7NNvJglTTr+f2Jn8LjT1gxWOSH
rlI1XmIH7zil3wQmqXGnSiuMfO82p0O4k/e0dRoVTU7w/N5Be0IqphFX/APMsPfPJGcwrlhothIM
Hg98ANpNpj+Y3ah+h5MwM4hTFaek9+gTj8MwGJlQiUjjaal56HBEiO1EHtAlVWh90g+VUe8Dxxj1
g2Xh6u4JA0PwuTPgXi/VpRovdkkRmgflgxsXGEsmuXu00T4SaZDNS6yIZ4nVthKx66PMxyXLo2vL
FccGzZZDzb6wY/ko1SsQ+NjVlWPYHeGWO3vblooTXlU343veCqofO1zvEUfJIzQxktQs5Y+oTqjn
eitMEH1MDJINEUTWNj7w630DUY/YcYjoQ51U6rBqIM8/km81qPjj2h8X4dU1iHTvi08YT6lJgfAh
1xjqRUUWtEWe1iDJvAz3C2khrvwQdNN++mwve/+FuSPuAx9BXSi772KlfbIeIkksl+v01ObYVi54
ZdiOqWyBTHur/7+Y2tgWaZircntMhxk9LX3+AAPzh3YRC+P08dHGk9zNc9VDabGFcHr6b4Y4ZGxm
KjOiq+vYr2XIZHj+hPMmA1srGVN0/0zIBgJLJNsPPcyjrkm0ab5usZ4T4RdNb5OXUp3VFikjS82m
I1WAqsQ1/5jMVDHPvjEyEenarvb43juV8q6xf8PGyGeOk7pmpe/y3Eu7JWMTIxg7vl2R6I6bNg+u
pWNl2/iLYbC4N7IIYci2jP/+a0Y4uMTUKX+uLVkIultn+DL9QLIhx2MThGiulhP8aQXCAKDEnZiZ
qKzvBexk0WVEb1xl9mUW5WRVJ9LW+LWiHArz/fH4BqGy0RSSe4hyTzq+mk86SB2yjVJB11SMWOi1
g2hWv1tKJ9p5SO8gZIfuzotDgtQXXK8HUzu/Ujv7wd+s8+7myDY8xNbuPJ6D2yVJ2QKmHUULAwjq
Ox1GVdRPLl60Gww3odc0/xAQdMCfl6hvvRXVY/vk3aZLiBdbcm8aRN8rxFpA4Um3zthEMSNEOYo2
0MjzXqZo0LDC+Mm/3UvbuFjqhdy045rC9iX1x8v4FZ1P6wqu+uPxl9Hn+P/Pb09zHSe/dtL0ouFh
2RtpwmRnj153V1bGqQ0htvxxf5aIQKVrp4W4Kn9Q+jKk09KNqMIQcfwIa1oxfuW9hyQ7luGVjbk9
ofyn0vbat1/QPL/1vnNAE/5cF6Rcnc4QFYx7jwKau9NHxqlydPPtHvoflESZvSeX+9ZAz4fn33eU
izvWJR6SAoVp5bi/cmgSHJ2XnzP4K2PxjGYe1nElv2lFDg/mXXtxefp1PAMUNdbgJrE/ooEchARW
tzg2X14Lah49zcUQTxfAt/3hX36U1th1A1hy7TwGMh7Sk+bqW26+/4dOlsMAYulD2xPNGM9EKuLz
W8rE0PajuKMJoClumZW71KZpCTeDxEvg8sNBPxQNxHawg5W3z7Eq0tuqV04oMJx1p2XqGcVKp0nM
y0IjAm5/rOqeTnmd15/O9XfbXQ9j5RA4FfPog8gwd2L/S6xJvA6u+bUpfQf9AexJx/HJTClf3o8u
TGNGTX+m1WQWQnLjAT7XPFMi6cO2NfzG4hUsVfcYKH3oGSiU/rQ0x8+FU6OyuKPmWLF8EpjhsCGJ
9iIjIgiDAjbDkI7KYZjsU9oCuk7Tr0jgZrBkb407yHxDoSHv8c9llEzlyxLVJAC6pSdnSZFilFnq
tV/vkNIufD6qfB/F9ocqPbA8SwuxabcKxWkLOLVxyzCfiaR3b+U/RpSXBtJzzMn2Z9qdYLjXYoxM
ZdC6N6ScQri2tRgiv4fy9dgzjNUghXauJ9VEU9z/zjfX2mw4iTejGQ0kstoHtCoBBufPO9t1UZdJ
X8DCNEobsEkayHcgarrAbNNLq+pOuWwe4wFRgom7eyH14HO5sc9WM9PoO597hbAZshsFiyGGeewa
rE4BusfluZp/xMgmRftPx3W5Oje5r2YBR7zoIIxH86yOGH711J/nrAJh+LJuLIz5vA8yaKV1K9EF
i9lElnRbCxR0s6Y8/Tu7qYwkp2e78AfBJUlTZ3ZMiYUkcsBBEWQfXsJ68qtN+e4eujstrz782Vzm
0GmceLTRgauyykrWDQl5q81dc7cs0hrcc/iyqE7vngWq1zfXjE0ZY6kSSnTkdcSqJiSaTjBAYjMf
2n8xzTAwrr+3p7kXRbaMe64Ayl9dDTeczxBgYhiVQWcsueQPPmhTk3R5AILO4g9iqsZXXeufsecZ
p5+txi8t0Ew64WdK0mxzf5tKZPbsv39V48fYsuR+E2o1iO+k3Bz4HF19zX/0qmcya0kxHGHF4rPy
bwT+vY2AtCRIbHpaw6qpp5PTTylkbcSpBVQq9qHKop5sXQaR61t5VyodbHxOyCY2L8cNKHUnGoH4
CRTu32K5QDP0qn2TVkTy8KZc6dy6oy7H198xKOcUZunRGSWC2y6EzNsyHX2n1Qx5AsXpqEhLaokJ
Ao4d+oW8deCfTjPNvR3U+gHs2uR6u2IsP5yIMSg1S7sWBAdkj/WIpp9kKv9UO2YSuKzgD4Bd+a2l
b2wZjUSDN2Uv7vAHg72ANvdWXeXlBEFtIY//VgBQ/nfFTtJhs/0akeSZlmq8UgZUdUtwliyxl1ni
R+z2rQdwN989KGEPjucujvjo9bqij7b+MK4MtL08JZ0avxsN1/IJzipe0T8UHFfy7KmKgQPbdz/B
N97uiWW5g3Ygvl/ySGRAPLirTPIZrOcja355edMzo6ZpA10Z4dDyBNuCiWTQLuOuMPGZIC/7TGgg
jdPNZfTbfKwSM6YDh2R6ApNsppjgHKb0OgjrN5QD+3I2vMPRdZEV5wx6FY8EDw+KJ6tRJ1zbSxo6
JRc/nXFy8alEo6iDlKkVrFq8ssps/WVv0DXo77lYQ9880z3HN+T3ZEQa6IO55e+laHz6EB1C3GOP
9N8dBAGEls+X+mFFVTAM7zRdqQgvbe3aZ/9tjndB0z9CI7mRK56fLpIwAqJa9ch+pnzhYn6OO9aL
jSWN8AZ+n2o1odtmlF0UsKuBovvFN+BTHOPRTC4sfb8slRenfPDGfvgvyIjli66P+N2jmcM5YAKZ
nixapKfFPfOuCtlzomwx3vpywGfY8haOMcCY2RPrKnnnntgScmJAhc60UO5wbt9i2QD7NGm182mi
ctD1/ervzXADDFZ+rWqa7bSK52KHLayd91j400CJkK+Ly2D9Js5K4WLHm8Pn8e2Q9ECWqSqYV6xi
uRhYAr+s1GwUsV+RGwdLUwdqG6wkkZ8w8wIhmcnEGUlZhDMh29NryX3LTXWgCZKQ2cUkRn254vwu
1ODsCAmjPk9rFsQNEsCfUXtoc9HPQlf2FuxslFfJA73AqaBLdkVGRC2f+RY2p4BTWy1qkOP2rM/i
MZyG1+kxaSS3IBsP+oZ/4BgPhvAuzf+pg5wJCx8MywcJ9Mn7FAF9o+8IqwWDDWbuQlgDbWBLDNUX
fdsyfk+TTw8F2UknHdnZHSvTywqYtljfkPNiG1rd0HL4GukyLOlGvDfdfat5FpYKPm0yLlLizfLv
Fc+/5rKbE8J36qXDitjnwBXO7hM3umjTYCQvcN38ehgY1dDDl8xsd60HGOf7co3l8bMkRNN++yrG
ouQBm8Se6ihtiIEswbx+v4XH/SVuYMA9IaLU3cK1RQVuD3U865aGQUdmbxulhatVjiDgCxil2ejO
AtLpng1F9pErIZc4C2bWoQx+LR6L9jRvqfABx8YUusWOLef+TIKgyM8jpBqPbgpkD4fdlunEXXYp
oW0bd0MGjXaV8v1xGFZmkdBZGSEydRcx5FFRwMaDR6fhZxeH09e7VCiOD8nHVw/7F0bLXdcVEF23
4reLzcvmLEnGmDg9/TesG7meOHSit94m7fr8m9fcSAqsSU4+nmD784IRu9hi+9wmrtZFLfJI5fun
Oz2hH+j72F7b8u5MXuL06TLWiuXjrM3h/0jsfI59Hld9lcK5Bc1ZGWaIA//T/wh7B7C6+m8RPmAe
OtUagwn4/EJ0yNJdRSCLOWcP6QeuKXnMTGwDP8MCnehy+7yA176kMfC2kHLBahoS+6uEQVSdD8IX
TB14hR9/Io5PES/8NZlurCx+3gwWA5vQofeHbM56UpEF2dM2r6YzK/OF7JmjKyctHk3/7eF5GpbZ
ZZVbFv3vv17oEPJNshZxc8QRnN/H9+BJ4jyelGC9YGofHYT33MM7GpLRWO1HQomH6XKOSxLOLNef
BNYy0MEwlQI4sLIR5WrFUXpKnyRQRkflZ7b0yTxVLJW1GD9N6Of55r7DBIGFuJaniBREtilDqYno
ULchhcYkqpmd0o26/W98QKc1EviVxxdie716Of1efWd08O0UAu6/oTLUqZdbLqYhgidgGP788LIK
fIidcg/J64CwaXsYFP1XMycAcRJaRrdFDqZBBWvZqBFjNUorT1zk/acrDf2qruCQQkcnSlPKXx1H
q12uOKEVTr5LCt+bAFV/xXrSH0NU71ei0MyNDGWvX8qzGC91UL6EdHr6AF045u96ddC4HxIXdckX
83zZEZjyy6X5j1kHOniTfJE00oX8gr1f4EluRO5TFXfd4gtYD3Xg5tszrbTU7UaPyIO0GzzmGiDQ
jiz7puQA2ZCBDtqYaRhmsrEEldIaRyi+GcYnaesIrcaMGB9n64lqrZpfVMED4adXtb4NuQ1vg1ZL
pTDKsKzWmSNCU4nj6kT+SVAIp6kOPxnxlF3ol8Gg4KLnhlU98QjA3lUEZqrJVc4X1nta3HuNAvlf
QWLTYQgLme9sEN56pcJGIfS0WJlCgzKiNiYBvi8IAwhF/8Yt0xtu3FX5d9hUQpUGBPfP2nJN67hk
ShN7B3ffmm9XX8HQFc4sGBswWJwMg7TTQyWPnXVcdigj9+0+0oxdxwhepy40xlLsnKzh1wR9d+dz
ZULW4mHZ/ildtwveLE9MOtQEu52XN6PXDcXwILN26lcqWrPU1aIhuMUhcFbTbaCCniLj5YFAvzlQ
U0FJxXUKjCMgOhmZvWaMkUpKc1FDEVYX1iJD54Ap4Q3I568ix3COECsoy54DHd42dGDaXgjdj6gm
0t9x7dq3CQ60pcswlt7ZEW0RuDTcdgMZLG9EQQEaXgQ3uzpRFqM9FZw+WxPchb8QdeHTc9i9dAr7
/IzHN+GedFsdf3Ypr9CBzw3j7sn1cHil4KcCkgf5/BvIjGKXsjgzcc4kOOBAhZZIR/tl6RLFw5Vc
IQQqV+4+fq1pLofYOwzMiDkSPLiH2xVQG7538YX+iF3RyYhRuD9LxgDfAf6x4gcBro04M0zKnxFX
LXrjgFOqc9NhwW1kzlwHHAiNqS2BTdwEvQaofF09I73TRXvlW4zp3OuwhaehHXiLhcA8PrETZiEg
o4g3hm+My6C6uzNUOre+PJxVE0bp5IQpfCdBg9uyuIvWVh9+F855KcUhQ6hTVhAbfGi9LUEWWcWP
Mpj9FrSEbV04jQkekz9f3PxzRhzqpBPwyre5xDsxGZnb8DyihNsQVKRcfVKnCQBCE6UwulEC8/3l
KG78y1oRcCshG2AsOHeYzk6t7oTWwyRpWvMvkyqZ0NhJIrt/LcDTbEOIJmgy/vxHwkxRZE2prP03
Wx2vaXIHT0ElrGaN+k1Bs5+ik6GykyipenTgLNqyLQRR/UBDgWAKVmbuQu44rfgzao0EAgEKicAP
CL/y4q0/3qGv9+Ua9XXieLIm/ceZSQeWgYnOd38tmTkNazsGTafT+65/e/K0exyyjaISGmwIDxXj
l/ioUidGgy4SqegX29xUMeAYiJ+g4Uzsbi8Br6CNAfylWHLnuGjBGEVpP9lsOCtHVs95J+F4t21j
J5NohDmxFHGFlK9iaXSjIeBYqYOZaKHIbqBRRAM0iY07hX+pkaBORYKJLMMoTOz7NsJgNjyuv67i
qQn5xoY/UpuJuq03E+x8iKt8rN58Jk19HWHTQ1WDKPealdtcQfIVR+GQZNG8YnF8G4pRKDFd/x/m
RxZWvaVOmt1xPUwcYYGrwNBCCXY7C2oxQdYWLcUs6TAT+MA7vVWtbBQllh898iXM3U80WdxjEXgs
JeAJWmgxZK4xaNOHuIu1wE8rmqaEwqa5j5ATDFjHqFa+zppt1ohrF+RlDwRXhfy1ssJtk/FuiTr8
B34wUl4UE60J9fjfSU8FzX8AyK8wGXpTlotWPqVS9qi3llbddoSq0zDY+aX5di90QLas0v+snMl5
lVyuJaXNc8lMeuZ5LBJJVco+Ea+IWbeFsVFz5G5WK6AiUJzwVMe1+KNHDafw/lUgbo0gr+du7NAt
7lPtKjfYpy2jbbg18ckYUaZqeyPM+roFRECY6QJh1bn/8Gw/Jot1pfuWntRYp6iyNvMeXZN1n9Rx
2w8jf039CtkTxnbV8vS48FMRDXIyB751k2ZE2BVUrOh/VqHj/gXLOGDTEvWWFT0PfDt4f0XJIFQ+
P8DBV0moIZdatyaFFSdnhqDfY/I3c3EjU9vau4z99n4hBNEHG96AIPEBreuLVAvuEs/sh1H2uh6t
9LN+qPk4hxpD/ZVBWdOvTggpman4ABMr+PpciH6AKkcetXH4dpV5li95lBaYDM7IAO07qPupZYWA
dlnsOnZnt0HA06+9hPpzyLbvaKteWonjl9dfBBdKTeCf3jv2kf0g+cs2Bwlyc62m5bOxw+pakwhv
zAc3NhhJ3UrFWcaJCqWiC4tEgydIgEqn4+kA2VnndDjbG8XXQjlYZjqcPmv10mZnwLwFKuxzyJAH
zswBOXbLJvGJOQQAy4BCQe/RIXQlCeWI8JuipOxOEN29PIrK4U+LR0puf3aW44HKKYEIuQVaf0cG
DddR4Annnsq4ZzdeXx7Gm3EG9U/KR2X3laHz8WfKZnajycgnSXK3XGrGf6Dc1j7+6XMIdGMNIdxO
vazxKsUBCdULMGmEinZeY3ZccSqZ6VUpA8GNleG9HoT5HK5TO3sgcVMfnr5Vm/EZ/Cl8x8AxQOy8
CYBo7DMmjW67Zns8zHC4B6AvcWoppsBbfqBnNJFswWrdK7/fgHBwxFGLvcXZg3YeyPXuk63dwq/w
X9ENl9hklK8JwomHCInevSVQu6oL06Z0E9BbrvIYk67OR3ponLF7h2mMPRH+2tbfJ57Do5xA4Svr
jYd9yKV5dECHoVRcIvcE+u8GHlMKrt7iiBMi3TKGJfY6WpqVyzjxq7KdFVVB693PKKS6xJHkBsrm
pB3HwApTuyPnTSI6lWAkT4gjZc2fo2CwNylm5/gvneKftFWtqydRkbh5J4zby73Xb0a9sGRL8uFi
nXBWP7ymk5m3jo4RlDnmzoq+nG1w3uTScFpaMyoRQqhob1QqcDgtvkizMA7mX/Po6Xkq9WYwMxez
q9FsSNILYRGOJW+kQ5EAJsOhdWiVqebbuh3tgU0VvXXN53RkwgSj9W3zxmgk4S35g7CsTdPJsoa7
DFpB5zNYy885IilsVSt4TDy2jpUVEbBtVv++LPWCvofW+1aMePCqWpPe+lEQofuoQk0kr2TcmMfN
4NYFDPaaJ6NhRT3Vy4grnJotvg1CWXKrktQOYSua7qXgqVlw5gJQuGQ4LNwwwCP/woj8cIQl+HlT
gV4iK/JQ901/cunuuuheewIzXOgEqCv/YxnwoKhxTeYjK8KvnVAZOHLnzBzG3udqw6sumkGWZByF
1+nKv/LN5ua2/5vppZsFGhlYyNCHx+KP2VFM/aFCxR3QRlPhZH2hVp86bfWNjgvS6wx8PsVsUa+r
enZtPCMx7aOiHRvnPemLQCXsUgrCljr9S32WznXlX1CkKOXyY46XebmVCWpE5yVyB3GT2PaNHj34
IJxXzj4DkaFHqkVpto18TYIAiy7GE2R+w5lPuWdpuK/Zj2F7sxWN0JjjjJxV8uuD0N37h4nymHxi
Lwzgry8djgOp7d82rZyiD/QJHLca+igXb4Loc0OCrnDE5kVpVQctS34y6dahw0HB0kNGeRzw0lMl
s1d5RppDLyOMrl5LGd+LCqmPWfkyeinDC8Mlad633zcxgB4MtL6hfEFFb6Xq28Zu8NNy5QcqLX/y
YhgXY4Wv0HsJ8wcBLIKTjn95AL6Y2a8hzVVRkhBNnTmYeBR1EaaIkWrB8hApBSL7Rm+nSAlHo3Rx
gH3YG5YCmTWL9QJ2eSNDlpGOiUQPD6XMatr+bJ/yghhwUWi7uCPl9SNnxebHeX56ALq5iycSifP9
l5JbwM5meGbpyGuHcrDp0bozRV8ucOH5CcGXZsnLnbPsBZJ1tRJ+x+l6Us0it8joV44aG5iL1P7P
rXgjqpoNUl7FqIZaWe9vU2/L1uW2+Zek6eoCCR5qrO24IXdPKwVgsr/piqcIqS2+pR8DfOXRswC9
xZbN5cNnlU/mQxp5IGjVBLjxK/TfuYNVuWOgpGI96U5c4PrWNJlyTDoMCVYPZg5L7fFqWAWaD0ye
siYMI2eKPKvUttSY8nNgHB24ny/OapkmQz2eygKVYhjknqDTY8rFAUHvFQE0uWUBN5kzYQ+zRoXR
LBfe65s4HRRVpI/5fBs1oLRErR1npY63ohG5z/kTNbKyzgtzdzRjWnH+O4vzMTJbcX1T4qeBDOFm
Ijk6YV8jRYzKiCBhlzr98potIm7ag28SSJXjNj7H/T0o5SiNv/CcNqGfLt0NiSsCkXtG4v/Jkr9h
oRx7WHVNlmd1Thi1NQroaiGPoVy9O42LgKbPpnJTIW6EmcdAcTztK8YvV2gcsjKxbOEjDN7AI2U5
U+HXJnpDh8fKzjbuA9I6tX5ahHg1zre1U4FicpKHlOXUCPYpd88ZoAeCSsCUIAJ8JFbqCRXZY4DC
8d6prRz+hlit4aIQa7lgNlI4/V6f178q9Ne7uioNVjwHumort6jHNMUW5vHi0MR0Ce/zDhd/Pgsc
qpvwQ1tMvmGfBDeivCwvxyYcKAXx3q8xhtQy/WECMffs6zMZi14zyRmuBq32JKskTdbWY/45W57G
UckefhjmLOrLOPc3j64DUv74Edk4nTy0C4vkrhUmdi/V6XLpEBat2JWbAr02JOP6O1Jv5ZzZTUap
B1xEZs+vOpDgWcEGXgR5OgS99UktFEd9pXx8NIIaj35/hrewBYLenB+8IvjKdWCYg8yZWkCaZLef
1SkY6mcbRg5w1P0tN2E6ixjX1Qv7hAvADQGWnUEri3JDH/x4hGgJqNDknixnwH8rDf7WfjtGGH9U
FPfKVMMAiVMW/RcJmJi3tTzzhWyEAhmCj8AKwP9X/Xm7He/ykqD52XhlIWJALRK3Ej9xgdA3XDo4
0eUVF8UR6+AUP4vF74WDVG/hBU2zEnxh/c86iWsEGOfmnQuS6sgCHQ8s2keWafVqwG5k429nK+7s
Fkvbm2ulJhPPGfUcX9jToWsDnwp1sB4jXf+BHr9H+mzHI90qrqJ/u8WzWaiIRWY6YrDCglz1FQ8E
H1dyvo+YFrl3Cqpac7Mx1LV9eyDGiRRkLaamFFaC5TmkEQt5Uj2/ulAeYuOwXitCFXXRPU53DtTt
84iqotKear9jlRELJadg5R+QkGojFo2MVIpLHYtn5vZOmiUCZUcPsOzFCeSruKGtvn8w97yEWSAm
yTQf5fC0XqPb4P05LfAuzfh/PYMV5osjiMV0h9iuRC6wZrFfuQ2V3w304yF7hUzAFS81fc3IW+dc
k8s+Jk4l+RrJJlET9b4vhjRKpAm1FJlafhDJT9Ao7V5yf/IJy4Yega3bEj8hOuz3v/Hx0iROBUxQ
npUaYIOi2m8R9GxNFD4QTI22JFmKHadrYUP/GHOnR/pZQ86svGFPioDggA/B+s3TQaEslWJY1o05
9MggdiWrAzBZ+pZG2PSO5KjJTu9GQLViHRqdWbzpFdISMp5SpfUOUPn2TZgFoizDWUJd5ouZlrrY
1XUOoyUK6gQu9lCqecI/gUvaqhMJMiovYazH36a2xnrcP3whgz1de5fzl+mHh1H9g8h8m9YD7rZD
xkpqSh1i0OiFNqJAGWar0MyAUaNGWxnsrfkc73ZR/0Rz2uiUu7XWi14rVsKZix02UCpDxc4iLRnQ
yRrwaWKDHZ46lB9gBe+fDojv5MwgkXlAqleFbh4qdxOl5yDYsS6l54czNe6GAtIeX4iTWKaDeDq5
Nk8ys/fVhf7+/tftk8Qj9A0Gk67ShClLi4dHIxk7u38aUtzvWAT8NKqTKmA9wStO0IjRMWXpsnDo
wGdZl9PjljDUa57emV1vtSKxU5fwj5bcjKH76oScDuZmnCcXESfoi7tLoeOg5JybaiBR+muzG3N6
7g4tdW671IV4rQiv7KX29a43hjZkikJhIi0FuyZqjRTkXUas9HCdpKCCHRsDz8/nAP3yrcDAQ3Li
1I2sZkLsVekPZW5Zp8JcV12+RcZ+6oYKevHy+uduNq3anTrF/jVSuFPufB9i4y6oY29r3KFYXY4F
FqHvNWc4dPRHiu33CEDAOMQccvgLZ9G98hM1VgsdZHXVHofCMEQMqG5pka3NdPc/sdRzb6myFpBr
VPHGWuhPov6R2/bn9HsdrtQeItEA1AOyawPmhr6KdL56JL4phTgj8yL4TSHpcTcLXfLU++tICm3s
AXR+HHxcHEkBs0e84kXgHGY6uowkx/20N6FmdDkWDTGoHir+4yLVDOSnXfeA/dTkH7Rgri8HECs9
HqY1mWrttCF9OyA4I7MSvTYtcIOYr9ew7EHcXo9SCmY9gKzc/LZRKlsUVj2D7/v+ZFnC5/OqHj1e
0HM7yP1x9ylxEQy1B3o27SDbQf7Zqwz12SnrNCjGECN9Z4VZntCTlXJHqROBmFDsxOl5Z8mcibv6
HE4rnn7mAE3Lo9YiLCNPgn8XvgwIvs1Rf+WJAThH3/PmHbshfI/SNA5zJ04yXosf7KXL39U9LAZs
vXoaHccmDeJ6RWMnn+Dgc/80YWkQ4URTn77jyTc/uTL4JwZ77gV4yftCVBWMpsWHM+YfwwEQyvMD
jWwdXaVId8YD/Ny5iPESMlhjoNodaCeZWImsU33rOJp5TPmfDhS9LwUuxOV1Q9Fztm9bL7I9wO7K
HVOMmOlXCQD+pMHP+yStBYjWCjWNecjCWFta7UadSvJh46lDhfoLH3CfksvAqDad739Dt/zYFI2L
WKBEYCOYFrmFwmOskFdMRgrkjFldYNF9dVq1AJevUlj+nL8X44qrliIRgfInRwV0rTApvgNaFtxq
+RRY4ia5g2uR1i+vPhwr00HoCBlzZ82AhKbERZncNyvQ5UNdD8YY37PiCcsWGhjzv+rtOwbUzi/I
xUrf/UIrPgaxlnGy2gQDSc/P+GH9KMuJBWW2Isme/MuVm8tUygHYD9bvar0sJ6eN5t2uaWDoeGPX
uR/OxCMEkG9oYO2gPFRN8VHE25JeOXimH//NtGTYRKnLoQMi+2dBolsugEJ/eUXHA7PLFWvCrW66
7rF/JIYdh87axAqGvFDLTI4O8fyplNHmfwtjSDq+VPshNruC8OEPr4DPKaoIloXVV2CC2jo6YFiN
gE8zaBCgVW19gttGfRQoPVGT7J6OfkGqpcWg/UHxl5tQ8k5jSHFg//k/nDpfQFd5cV+c/UyR5CZv
5ExSEZlPLDQUTCzrhfBLUwzUp3t8Cr5R7I6eDrAt/gp88Nimxu6uKYzxMyHKrAQLLqrzYwix8dLU
o7/UQTlEhIZ/pgJnSRK/tZU8zZFS6UeAlZkHmB5qKpnMc0y8+9tAYGbFvDcmGmseYDalWkGPZ4xl
Fq6vvFOZfA6nYZZ3FEeYnAoo3oZ81FKglXeiehkfOElQQjvyt5vDRkQUY/Tg3Qb1cY3e/WWTC8Ks
hD106L7nC4sAiissdJ3jzg9fG+1CjmiWl9xIx8fofAXC0JZ2ECljCNl4YYN7NAiE4Qpl7tgV+oOE
1v+MWzzAtI62o4kIofjLyaYLyL2w06VAALhAuXknAm7SVmEIxS7ht6Ag/MyiGx1/xLcWo7Gwx4yz
+23/0Nr+avTuk6iNCEyNWhPABwwu+AqL5rNruwj7N8U76MbGuOFriIJihu769tEZVpYonrW0GQHu
qMYdwGO8Uf9yH0jlj5aBzCKmf5HCBxVk34lBFTUFHWu8hvCKmNDc/yHaODI5gfLNFNz2Ax13wE8d
x+qzrSO3pC59LO7sn+YidQlrbi2PAkfZNsqc2ype9AQD3VoFqL0Xr5w28RIeN8tkBqgTbQPeCIAJ
mYZp6/uhBweJYCAgllQt/42N+blRTOAmH1Jd8Jv57uynZQSMpb19gWX5x40i8Laj0QzfYmiylmri
syrQDYX/QrpCg7RZA8uLSsc+1J7dztdvcSQAeruLdC+nWOSzg7NqA66e1XC6xttR7r+uMrTq9s6e
tDg6G9NcXM84cEtm+m9QMSvZ42HW8St8cZbqFl7+kzej8AZpgwt9pB26wXYH0rv8SpPcd3Yj+XIp
tLBszihTr1PTO+e0iDizP/Lml3AQ9pNrgODFRlUKF/pJG27VGO/y3CVnthEtCIIcrclqlc6E3Ssc
Fg/98g45LMBXvm3tDpiFI5W5TU4caSuQXtTX110GKFtPmqyDk0jweNmVnLZlbiaD1mechyrvt6Sj
W9LvDgG6k/ulvjrkYFHoPz1v3D5t84qyTkjQgmImMbItj1v4xdJY7Tk/FmryB2Vmq4nzWDWAPkqG
zAtf1SMgVhD9oy9uP1srtPPA1uzJMR3CwHVJrrIBa0stBa+aMZCCJTQpQ4hmuB7Sm4H7oFbYFbfN
jC/8IluLeiw8V386fOrPptoVlytgvmrFG5DJE3myptx6szD/1w7XYeRJboGMplPMEvEaVsNwBu6T
m2Vs5/N+nSQsUSCEWIO7kRcsADpIcCzKAZvPN5ZBTWw0mWsR/4FrQb/DM1evGY4Kr45IXWp6COMP
rY1coEEw+/7A+zIW8xp8E9Jhfoj9LI4TfDJ1IQ1VnHRvvtHHy4j8XDUWzc/SM566lks7QemMHorG
gJaVttXEIfw26JS3hWopREnTEiXfu8kpbGhFlZhGbws23/n/g9/ZXfISu9rZVpGBoWLmE+RKO/Yj
mQQXnl9grr5I+Y/8Ke9Iouhjeji7ZlRCxjqJJnNh0Sei7/PE3dIMXhbqQtL3uKnodpdY61iKNrrR
R7Ph3AMRPXOwe1ICodw7RbvzAPRcf9aW+L0WzFmxSua7/Ts7zqcYr0AlUeFmHnvyBrm77GOmoVvh
l05LT09+F8ZJgbjTiJbqsJ0CS469Jti0UVQiGt5RzhrLIBxuOHsQx2egCBzRDpjSjfRN2lwZ8Jd3
3lKVmRUnReTfL98RuXjRH7K73C7M1l7rirgkgxrrgmF/TCn8z735XcZgxD2TW6l1VVABLgS/w3yH
9Y7pn8NOzrFpBQgcwxkEYfohu4OlgRka838Rr2md4RGCHSfK+BCz0AQyX7bAslKY8T5f0m966pr6
JOJI2xVBaMLv1dRrwA7dBvB89TvXtC44eiTW3Q5ObJpuQN0TgbgO4+Bg1XuLzkaVPS9VHyz3XJgR
Lx8DWw7EvAPOdrPzuJ883PrZfZvBZPa/z5bIfMCCF/kqb6Lt3q3Y+Og+FYAlaaTbEQNyIxiwxyFC
HFMl5UehY+5A2Dx9w1tYHQlRaJuaQm7XpKy5Hgxp4rrGM/AcBlVfTrKEGB2dmoYFNthYLl7xc29B
U3iQKcVxmNcl3NTxA7h2gjoxrMLXRkkWaEM2KieT2VrVUCY0s7bEAxU9SysyqASTCew5Oh3EplBl
pHX96CuMg9rC0P3kSvHZ8XDKrlKiGPc/KtZmt9HvzRcrXBL6f1I5FmIiKyYwCuJAq61zxhjLYdoJ
EiQp7RekE3ChUrvQEoZkcSL1fTjrbYaw7KyofMX3C7urKLbEkfT+7Sc/CWxbnAxhBlfSjwhZtH3Y
azeVcX9wmIEsWo/KIdd3hMfExD1hWrlS20STKHRMnIuUefxKYTjjSK7tqSf80NJGMOlC56Pfwr2L
Nr6fI9b0OMJWh/0ZeP210MDdeRIMParREi1vTLFTE/3ICeYT01PKqcpGGxaZ88G3OJ82Tt1HCbip
9goWKQ7RDfdrAJG+sXuarzD3WOaMCSyF+57fiHmS9jSN4dWktV75H/4Vd5Vjt2h+C5TtSOSynTsq
fqB9wRQofcx9FCdMffxoP9fQ+xz7gEyHZxEzB/uYH+aOiRCroKPqqg4KZZcpfIw80O/ZV4v12WiD
coKTnHgd+hbcQO9LxDfFolNZtbUtX2qKdy5B3oFPlYHgQF7k/6TK8y1Cd7wonP1RTQ8iX51moDEc
0JUENRfPZ2TlrnJY+5TTJp76sMbxR6je3hFrBWVpPVxndlQ/0Z0nKt4UF6nKpwb1S6+jYpFUVhE2
IP3HkbEysqSO3uE1jTO579R+K4zeHBvv9dbMmmYe37rcbmMEX7p65wo6yd8bES3NCVF2v59uiQTz
GoEExvi+5FFwvQaz0KHEyWmPUsBS11pzBLpFUYQPkltTdcQKBtVMTqDRrnT4wk2BYno5YLutNJAv
YIHKBuHqwL07T2q+JoK0twnKDQwk43G1E5sNQx3Koe0HNYbglL2Rnu7COQAhhmrsPZGnAkfUucEN
mbdv0eEjp3j/8Xde3bD7v1VAo5Ge9P1oXGJ8Nm8dZtpU53dSqd0+QDeL1AuplTaOS1wnwP81Wqbf
sSQwKw8U6ezyj5U39zoyjMeMKtLxg2n5+FCzftGGjchAUOevo4w/79rFzWueaGglJ4+KoWZIFPvr
Hwu2GZOCzqJX/dEXYsmd+LXVUPMccSnIaW2eM4HQYYCZCV8hdqk/iKyqix9gz/GyJ1fUaN9pvqS7
ch3CoRKJHHvhhknvbQEdbz7d+Wro8pW5cetJOqVR3+XMutsGlozse48MT+9Fstsc51B7z7eXu3mV
faZdY5sE7WRQ4Jf3f8FthXIdR1evMkFvLnBZbvO9boZHL7jZ3PB5efOqHhkkKg1i603S/69Ym6Ui
uf3HVvbJgc0Hn54dYMWBXfrr5BwjGLaUnVZeV7I1sj1YRds+iDjWJAO60upvYFvi3UvndUxTRtu4
7/TfD1KFnBl8k9Zd7b48T+QE4JYGjOKQxLnJCZk5fNCNGXpyxzhUnZl1+/wOTYPTj/Ir0dmzlcpL
stU4Tjj7RIXsb/ZVH1To8jsI9XApwJL5tLdyrOljdIF3yogCRGRlZzJWydTrEZhLVtHPeI+MVrre
24/qcQgAx7ctPYFzhxHCyAzAgwT1v2xpJ3ngtSTTeNivsCGrasgzlXHWB5bPE86nPxmqIx9WLe4n
AuuFW547bh9qDYHCognAsG+yB4uiOfqFYhPklmZateFK9RQN/tsNggFpPfz40YOVdXep0fhRJc1J
dsMXbQR5NDgVrTF7fnAHuEZRL4pNikBfTX8sfrVQoYs/PbiMW3I2b6ZufItP6QJ3OkqWSMWKCa6v
R1nFXw5TfcmNqDI0+pCCyzVcwcqph6DIt2NBMQAAbUt1xtNLCsVGP2YXcRireMB1VtWwO3Y2mn43
633cq0PbqyWrnGiZkH+JYNNKdY+9ZlvrGm0xJC+nmaIT+FCKv5NyfsIH99M7y8FAdcm0GfyqIL7q
rT7NuK8JbzfKQ6FWMxgQOFls8pO2XICIhNU6b+3QDa9lw+Yw5qmifK6s5v22kZmCXDLrg4Qk8a0L
dDzhh6KzYan2rGBB+CKzKGTyezkjYqO56aJ2LSAkeXkCey9pIVsuD1gsbE2h5ILGpvb5me+5ZkRC
NU4I368Zc1Uq35Et456spz2pmNXjq2cJoWURfAiVt5/I0qej8qIZ2hc7aoplZHRTLa2fSRgBh8Hs
9bBpqUnmjLDJS80y/qZaRv04/ZB9aMwmDRDDzucUZo7NoUVrsq40sbBLdl/bxL58zNowWT3xIoa/
MKEeplTrHmAuOyqbQkNc4SqbVodEfoWl6Edrn+trnnSYB130bPqpsF9NtSi/Aa8mCHkpLz5zTEq/
hb3AtvPUgNm4g8rSsp9oqo+LP+KnqZWuugBcWbzyisY+95RAvQS56u7Uyk89CM2o7rGisOs4j5Ar
86FBy7+YyWE3yvpy3K8Vt8/s8a6Js+ZMv9EbU/xRoNhGmPn7dTCGrZQsw+kv29L0MMxOVm66VK0V
XT9pjefQ/Ukej0+N8bz1sOSeMXEtu7q1WwkeZ+Jd9QvqvYnYms4V+Lq+qyC8E5fl/kBkDXEp8m2h
9HikSzIF49ivIb2mbsabMQYB2N7rO1VkEZKFEuRnbP4zF426JEYi3qr/dpUd/EtZ0Rki9sNsXGNh
gxrrAGNeXRAMD4LRqjsTEhRmCvNlWktruiLSihUO8mYT+sZyofRsxj+wHNDIJacNUiPKTh1tYpBF
u2bt5qs5TgV0kx0lafJ8wtKtjB4yp3+VIVgkEMICqeUaDmAs1KMIU22v6qp0ah/wNaJN0fkQwZZD
QlgDCG8/O0uJ6StiDeD31GXrp6v3bJnZ60o7hcguZdDdQGUeSjh+oh5ZAfa4j0o5WeWCAHe1f+Bp
X/0sYo+OdXI4c8nwlia0FbjKbZi3/PCbcNXZl/cznQbTrLAZbH+uf7xgZM0udqYuXDoysO1b8Qlu
72orSVgJuAsdNLrwAC51vKZDt13z4ba0ikN9bUAIFYkowcpoULt7DCjHCzg6FcEFFQN1fa8qjQZe
r7f1kk3jRuZdDAjLuVzm8G2wz0Onu+KDiAJjFk2FFr/QVbD46N9Ysj201ElBGrswjYWJvzoLyCG+
p673eOIGQoZSy2dMbK9rTVomVqY2uIsJtE2XTUfXxS+5vgfDA0S2seXgpWA4JzLGcy4VSySutkcj
x/fefgdMGcO5lP03Qf5gE3RDlnXUWwveELtVT1hRckOfFHrDxh7qKaDwqk4bcje7xBhWmELODZIP
M1+AeG7A3awdL0ozPd14VIv8MlbhIveDOyGipe7K3bSQDlQs4i9uBM4wgkC4+gjAfpKI1puAM+Yt
eu80beIwLkdr1OoiApGAwBiRuNxktPn2S6aHf9eGdA5/QMxlvnjE2tsHgTjoVzwHDljaLnSV2ZOt
er4TeFm/dTuN4UC6LyMPIDXqvZ5u76Vx909mb1v202zy0FAUAv++WYfAmcLNIajgxr/DH+Ci3PaS
8Fqs+mhjrFaFe5lkWhPL7jMr0zg+ir4wOeX9C+s35yZmyarqy24+8qVJe4kOCpNlY47+AKvhdiR5
eGsMqHp2tZsHIZmjsfoOpORKbmmau3XVn9B07zeEJzK/JC4MRX6hqhyRvCOcKWilHxu9GeM+WTUQ
jkwokiRch+8+qDjo8BIOO2IknSU2Bx3BT33nNQuAr8WdHMrnQdbcBlveEq6ajAK6gWVb9CnlR3qh
TRdlYpBR8+7EIgTSZQgDSbTPS4JnmFgAno1Xi8giQD2i52H+bbCQLKyrkPi7dD4vJbRNmByqmxNF
ZlrWAOUcAouanqDqvM8jEZtXfPfLq5TRBn23b4yVHI6Qb09gDKyAfgAE2A7fmISM79B9ITenlJcW
QmGlMX99w81h87BcHrXi9/bx73aAqetPSJg8iRJfbod0i2IsWKuewVPk99ubZXcfVwJVn0r6IiaR
aiRqLTPI3ZqybJPEgC3U78oct07Fbu8BWRQK2PfNGpHb5dkyYfKO/6F9zDGbKr0rPAfXQwlRC5xc
3vvK+4F4iJBHplsrd4oj08qe+pA/ykHn8jXY+UYqF/AfXYaYff4NgT6ENDEPOQZmj74ahKR2C3iK
D5aiTKuSch6CK0PK7sgsB+VzAN/R/kpvtSP/ZeBrUbLpuz8trOKhY899cQFuJZAJG6vuA7CrCrjK
aBT4ALEkQs+xRO9O36Xh6qiuTjw2CwzpYSP7ZeB6QyFinLuaLgtwfxWr3l7E+UqgEVHj3bNv+2al
IyDU0MStjwJ0Ppp/0ArY7aYqalaDqQiUFhfDXpm8ghMGX8+d9O/eOlnKXOepGe35Gm0COOi3B5ck
hBjbkuSCs6dm7VJeRMS9LfNabSLvs8eEPXPqAQNVc3aZ8raCfTwXXbAnujWcvQi3mc/3ei+LMn6Y
YCF9yE3Q/QsTh9t5WohQAw0wN8uQgSmQiYVO3nW7rAFG/LWiWOOjMKHgMDlfq4+Lr/lBjn+CuYM7
RGa5np0TZdCFhKnQ5HJi2NbXUEl3j+VMT1eJeqTnTyjILYvzbNee1Grft2iUK9+MBEVLdALQaTHb
rs1r5uO6xEM2yZav9F5T70CaZ+YcS8BJslYQsBitqpVAOqymwjw0Ml994EXkqstb72oDYVKmxc0K
aIkRE0Bnoewvx+CFJkXVVQBECyMp01w+5vqJ2AF3lsVXl2mr5SGQeenm9pCOzo6gbPO4Xi8GUjfU
XxKvrd/XPc7khQArEtgA/CqTkpc+YGR62OJ1UXzdgnJGSyk4tQVqCMkggPk58g5xdq/MUYFgahAK
b0Y8VmrWPIfIytAeAULsZrqrBtM1+kSmGnF1Cm7r9Lt6mLB1CSyiRim9hCFm5c/J8PCGDPVrUs5E
4uycIk6lozDZ5RiBtgPRMTY5XE1mZSjj9/cNtc57iAKCJ45BDYBvNVz2HUqK8nVfsm/QMa6MrfSY
8otZ5ucS4SJhM2YFwXYKWr5MDPTslN82Ud364lLii1+dxQQ/GBcMubW98LMyWUJGg3Z10YqYVsnr
0jV08LDHCexmCVlXNHXFOl6PxVBH6g4KSykQWYuEt1AQT1wro11QdgMFett62XPPM0iyk9f0hGXK
JeIEcvneNuhXxybQhf7U+cVr+p0CC7xiu0DKH8GRNRKokkm5PUv7xNJkTp8qtYMvhKTaFeHgzaEY
2HIRyp+xv5ptvsqNcvbL5APN0u8kr4XuGBmL1ukpbzmgm6/V8nPfILZUZTQmG0H5xpco78vWbTfS
I5siiww64kXRYrBDw+0tj8Qt1dDjHICQDN0TFzH9TlQL0luZJdbZNBOlrsAl7ehjpXzAyTU95leN
acOJ8QC2EH/U1sjzQQFfX0rh7pakxsiCRokPz4rcWvXqD2xQoUiCcvAntyHOOqu7mRkwQSm4nqSN
DlJ4PhcFstbFcpMfmlaINlqEprrifcqs3XktkJE3I5LIVpNTLX6uYS8UewsVZrQ6p5MtWIrfN+4t
KlQ65hYr70zHZL7KiMNjQ4wBgM1xzeuWeD7dfK38LjRSfnX+rNIdCTBYbU/rXbhyFWfdDaKUQUKC
0p1R9le5nS0tQ/40ToPPSr983wBf7WlvN7jc8TI/fn0xAdnoMMBACEu4m1098ZNVnSEz/P8+JWeq
k3hILthjenC2J3pObEJ6muhmZU79TzHyjEfjDBX/tVUNzhbww2GBElMAujRRVUlIOjq/NFRcvc4n
UQitqYb+D+weA2M8pF6dUkeQPfSdJGzx7/puilhdmTDxHv/aj6NGyNfNYL2Xfmp0OzX3cwW8F7lK
UsSBZXELWGOgcDwKEj9733GLFasZFChVLsn+7oFyShtonQ5Rn5sIJp8Jdj5t6P4s0Zqcs/luAMJ4
fCOWuNFvoqb3tFJ8QG4srSUAjUs7myh/DibmVSeNik3vpZZ1r2SLh8GB+te/kJxSONm8L1/6mALk
pFgWUCOsTO+ohEZB+HWe5XI+VVqxz0X8HfUmqJhRPuWsY4IMBTtEBMbSVvVblUGNjpz6KtKKjoMV
ahhJzWF7YyB6VjAZy7eJPiZvoI+5rjePZ6sE3dj6j9uCf9ik/9FFDBAh6viQXduGkdyeoxpxe4Yr
EqUjSANV6FeN6YK5hTVe1W3GD5RzBkoJDzwtMSkLAqNJplgNWBy4XAl0dJIvAwKXRJ75Gd3m/et+
bopBF2KnhnASCVvdYWgnL2G6c4dYqYcKW4qgcmhIwgNEMVyLnWwRDAQ8bDNzmqEYVfEO14AxYE3s
hWeH4ZmS+rJB7NaOBRHboExteEwfosF54OxI0dwzGynxQqnJaIcvWkbSDssD/GIEyi8bnA10kvbp
SAQ+EY4vgfTqSXp9P2tervJiE46iprYkQBCpOb+uqBfVNUlMu5d1xYBpWyrqBzXIVTXudnvSIWfD
P1A/OMkZPGk2w26RZXzzza9s+w5OxAQSDoZKvYCNHu6C5g+/OPtidtGpG+WKv+yh/gaIK7FxiJy8
nMnJivOk+tK0LiCHlXtUQRsXx5DE9mflucsLIbGV/cXktuPApilB7OwkclVbD+RkDLEz3vKc3xBZ
fKgYX/m0oXWCTiVp3b4+jXYJ8li5UFRqI+sVs6nuVZWJv7b1L+MwJ+6nTiVUWPXtWphLq1nljtiw
OfBhdszZnQQ7MoONX8/0/hufq+pG6A3p6uyfLTrPM28iLQM5D8xOfMKwcI+m4dZNhC4M8fENpVvK
hlZaWby0C2GC+1NSzThgtFF7RYEUlJiaE7XoAcFbsYoiMhXj6aX3IAA/9MHVqDs6r7RSf5+VBx7D
deanyOHMaskp3ZjRnJj14Ghw/03Hns4YZJWESNhxFfTLmtQ2Gh3LlMyS6TAJC+T6G+TbD9DU9tYB
7fp52EN0N1KoRCGyUtFeqAAkkRnx7DYqBpBJc7IYVJanXUP0ZWNZSpdDZxse2Vf5uN9d3tzZnRNg
NY+tzEcF5Zrc4aS0tfXiwjMgBD0U9s8N1vtXVlVlpod22GmBrG1Z1Ia4L9wKf4yFYF8KDXGKwP1p
6lifHj76iu0aXFvGCDTWV5Z1/aSI/2iVkV3oAU5Z8N+cEe32ziZKQTqrO2uWc53k2W1b79j6rig+
jPUlmxaRDjyZaHN8aYcO1vuE0aBzkMYgMBg3cfLXrmyBBcafSj+UKr58KfhrjiEVbdhTVXKBf0ru
Vxi8fYMFvY9ZXTfZ3CFVpxJi9QLK5978wrEisYR8mcS1hZtlp0llAiOLYkdDOhnM3hq7+n4bSuOJ
JwUdOp8goFZy7FkIoy6cYMNyAnNY8vZLAKcA/pHBd7dWDLn16I9j6Raml8Ws/0mnB1ojelJNdKIn
ZB6j7kW180bTEioUQrx4BAH47x6b8O0umSPztWivJQs/LzPRT7BgufYLSpZmPjdcqvq7+PYnG/yJ
0FbWKEnDWXYTROHqUc7SYbeEosWEo5JbUccltiQN/hZssUATfU3ZKllep8ASxUx6JrTBVeiPDWlW
QndfgA07+C5rzQR3Y0Aevjo/o0D6CppST3EiA7Ddc8r+KM5JImbVslB1AsfLM23RzSGDiQXPGpa7
wefARrHHYra/BXcNJvMxoXGntgKFT3pMNYpWXC3GDK24pMVxFnmfpypIIjiT9famnz+dvgjNWwsn
XnBP+090T83xDgsiyjUuhoIYJ1l8nfkH02ZBqQSYUDteW/mclKKJKa8kAnCwHeqy7fZw4U9gw+pI
HwAyCO+pQZvVJK6wvDYs7IiXJnbnPD2Su1cA5k5wDTaseooRVMTDr9danFxI5iMz6hq8MkMd9dys
UNSnwDo9JDjnrEC14D9oUuJ4vvrMydG/AT7/hTDt2fKVOcPy59smp0Gd6IVWrmzyrbWFUosZUN0b
bYFnLrPOKJXl9nXcM3jqfQKogyZFl1GO5Nl1zVcFE8GYnq7dIElALuUZ3B3zvAsyN+vrHLfKbNWC
47x4cymV0OhwxMVG9ErNKf/ppYqouBYFhYlieRxmVAbEAexRAJbsPCLkkTPJTAjSGHD9THMm9dNP
XHxRDdTbI8jZhyYl4G95blFA+aOn/UfNqGnVj3kn8QuKWL2rcbAayCVqY14aXTN4SB6M4wI96d/r
zvG/EkPywh/lta6jSlPQqTskwtG4rNIaE7cPqt0BXNrY+K6X5DmeaoJP7uYI5bDm8kXOb9sO3Mp4
4HVHqpQsJBWJ3ji7848rnWeIxhsBXotFVPMkr2gqHVx5JwwqveVd8iEoiuk6Ij7KfSYYZRR1hXlz
/ZsBKPo9oQfLiIap/Ye1e20CsvxfEB6GQqEOdAurd/0ZEvknSYPBzrt7ikUuxlqek3J0/4VBdlvz
9dy1eSkta/4vqqYEdhOKN8ur4Rkh9IlBNJbrGmbYl0nz32z8qkoPnCysycK21fkvFrt6Hd5HcI7S
EzEGdVVRzGEqABId/QCqe99pyBH4WpTxvVGZkFOR9hfYaUXM2zNm40P05iED49ao6rr8fwWwxRnP
sMuzMByusCWpIABXgKA8lp9KLTxTk9qrOHJDvML/tO56Aqc3S+yckFe6pBQgQK0zbz/0zNtDPS5L
DMS6TtRvHFMQ53/B75/WHwP50MLlkm5RaTgpjmbLQZtEOxgs8Z6U7IqjP+UYyTHBJyMe0hDlAFIE
bSyIn+Hp41VtGBY6bSIiGRiBFk8QRVD25+2dK3/DzTcXJDvobC4/SuKPDeciYMgD4+19Jw6ScKn0
PD27uJulJVsjci30OsKGxuc21upCqpsMxxyDejNqcWDmMSLRfLmWD/3X/9QLbSV4Q/xNLbG2Zx+g
j0S0RxZ2bsMi4Sylc84wUUmmDMwatYB+G9Ndm+GmiSR43zNEYl1D1ANISCLkxyx2lXHhnvTEqOk1
3qBRANBpcGJ8HQ3ozlFtjiMxHL0pRkCGy5exeZqCJUF2uwkWmnzHnuHNfr4LVv/Gtt7nW2z1qBGP
o1M/CftYsVSPRJMCofCOJLobMwc9nXAWIzh9ASHw+GSLq7cONDY9LFYPfso/YIbwdq4Ww5w1oy7d
b8j36wZMnjDyvzYdZLusfLjABOZFWCsmyg3uPWovM+nEymRvWyHv4MTdjscwhfxM1LWfNct5gav/
uDzj+tFusQCYuzXLhwG/HhtqptFzLrujgk3t33pyomNnW4/pLmN4nBif2WFtCCakx1uAGzw33KW3
/toxoOK39i/FuagX6bCmGbAaz1Qq3sd96x4/W1oDdj2EUDmzrcynMCNlm9zXr5azNTFStyS8Qodt
DHJfa/j5KilRZ4B+0cSzTaZ4uaSzuGdZG0HvrqgipXS6+JMd/Jzh5qBVhyCJAv5687PkOkB0sV3x
X/bNpwIOHE4t+CeXusOrzrViJ5ccl34iwvIF9lYilYUX55tupjhv759ivBsbdwxKQbYusHP27/KC
Idc0c3/moqCVTb6rCESL4ao6i9y3/Nkg/CpDsQV50XK/5SyBL1CzyBAZlqwj70EozmVrZYeqhX9H
dBrOOx0Hk8qLsd+f60h6/SaB7/VGrMIajKgWYORL2uWvw7VUbNg2wvqMOmRi0G6EqBa3uFc+Hr7s
g1GBX8+LYdetRXFD0JXy1JSX+bcO+OewTf1iZrwuAsP91gD2KwfZc6RJgtBS7xFdeco6ePv55T5v
pGFD81jD6662QZdwo6Gz2Tt2cgDNV2dz9fiDrh8SSonO5UMDPJAeYq16dnXoeUIf47HtmcXgVbkb
EWK694BDhub4hAuokHsZW606Dnvjo48iz4YFka+/yGmJFm56xLw/K0WQsU28e52bcsYRILvv0oWF
dwhztCZ8JbtqpdZL8Wzs5HSSLZCCrsGviUwZ3iryAPL3Y7a5Cd+0tVOfM/sABvfWzWeDiI9+JW17
mSc85Jcm0KZfHu2ImBcCLF9C31rNxCqzo968W0ACGUupZ70o7fhDOxOMQYqnSHzywBMcQR3u/huC
CAWlnhFQhhsZpxkMOm3D1R+EhyHwDmNu4TUh3ZsANso4BBPmzvtlQy7RW6MtqnOel/pWNkBomyVl
/kY5BhBw0vBpaNvX+eAvZ8xJ5yVBGk91CQVVUSTaURU94P4KfP0g1ANZRxqHWvZ3zPm9OFDQbniT
gWQo4AOoh2B+wHm/8DswlQt0VGkzsMjN8AIiFTnwowSGUixWq5dvpH9SBamIsTkyFQzxQR3sp3WU
BcEVvOur7yCzk5JCpgoiWAH2D4+Iilutxnx20ISLS+Rqq43gas+pF1si8mCfPhSkz16dOmJTPELC
ePj66FxuBZ4Q0CTTmrwgxu8I+yd4oETT4/iwzs/FXSrU6NHZ8FMPeezrV9iFztKgVSLdSFp5H8bM
GR/F2y4CGoJ3O9jPpyQ5UZ7+OylGFdRAFzGcSMZacrn40S5SjmWQ/rOGzHprjlGGeYLb32OkjO58
mVsYEtxwTgBfM7YVgNXawjvrRPtsHVY/JqJJOcvxzQgauKrUZm6rxgBZqZRliHD1LaceJ1BNnLol
IfH0GY/pQnCuJd3YGcnr3iAxPL+hkV6jPLAUcKQW3VPuRCSaMVCTS1lS5Jg8VKnfkgeQV5YWdM5k
HA444chD3Lcs+zbddh1Cx81Dg6x/O3yY98jMTHW1ZIxxQR/bkBQiuW419ytGW71In1LzJ9tcY5Xf
5L5VeZMEqSrTpaXCE+RV8h5+C2qbS94lErZZU9CHVp11zzwIWi2eCRl5WDF8HxQ9IR4E62j74qP4
cZ7JnY0hoAulvxPP8weIX11hVjyrUgttl8N/EuJXF6GeTwtQGSLKmwU3u02FUuAyWElVFPjzfq0q
kNGGUFrQd1ASGtNipg/7LELfIYxbIgzYJH1vAP59kf13wpVsIF90ERufqw6dnPGq21qN55+5J1LF
Ej+PlMPnzTFnKAl8VdrevtxuWNgsA+Ju4zMxTsTmM5m2RnTCOYpeYPCPGDXgFfim2MPs46glCllU
5GE2e/VxJzuIJpkUk71C9U265j5/JbXNQAyLitJC0Jfo9YvWqdBSJXLZnw4FXmQLKY5bLHJj43pY
xJEBSciPhCPpNMinxFYHVlohSb6QOk18npYOenVmsSzE4pHcy3LHKGsGUANu8p1SFfANeS9F4SIl
YHVNO2/oDNZ8M4WLEfKI7w5sxhNazoN3xDUbn8nItpNry//V9bvqZuJbH8y4j+ltBEH1yXKPEiZg
MA/GAdBl4WqKaUVBGPukzt0QgD0xg4A+M2V3pQML0Zgd6FOAQuTr/mRLFUd+dch1Q++/M9/35+l1
TN+a8FDSkYcv2MR+u9O1M2iJe8AeooLIEgPnei/3QGpCch+zWWOLQPtWv9U8ddllCDQ4ED9MhaJG
yqHahibno5f9/b77om/L3BB8BEp2klgmqEGzbtzQGo1CGS0FovA3ohmgOc6bnySoCN3HfsgcveVW
D6vBD0wKuo/Zsb8EM6IzjVA7EKTpI2A5mTrV4G/P4WtvhUFhl97u7G+2ubmqhzoqPZi1FBCDir0p
71rkUYGXkM87X+y528nV9y46R1ILx1VfcClk1g0Fiu0XcLLo91oCnVHAmOZL/fYU5f3B33pMZSuz
kFxLoIhmtXjgqgcSw4Hhsgwe1z8K6QuUqMoTepPyKl9PX8yEwX3fy4I6Ff+lhVtTF1dHoo582vT/
QpGsgooGlu5hHuOkF9eG0XbAPSnsIRruwvQjr/uXrTJtjs7IvovIHdSLZPbJ3O+oAsXw8/Le7NEX
yGOgkNxhBcnNmEIrC6MaWTYD3ENyCRne4F6+pGEugWTAc/dEEZ5bNTaU2aGFl10Rbg9v3MYD5ms4
Iq8GICjvmMfckIekB5C7Alaboovy6ZPqZLqzHHNjviMO4QBDOHkq9duNFkrTE+qOr3s2kKu+dsDF
aIWpgD+s7VTPv1liztAeBvvfJ6t5HzpBqigZw2qPg14DudzxBOon4y46ZOGkb3TyE0a22dbw8osR
88CIpnNkmIWDLm9+pdcW2ItT4o3FuZ3t2zG3p4w65EOz1aHDQWvjyilG7EnWlPZw0K6dSxzm0qkh
ie/LcWzyRv6EAwUy7tVWoatdLv8iRIw0ZtrZKEIRdc/plprh999bg0DPDnmUVCUGZxYc9BTmKEw1
+l5Z8e4RUkpHt24+ZHpmJPMFRfnWxU8j9MqWjPlM89mrga68509m1bexEfWXwOMK3JUPyMlPouc8
fTRAkpLjr0u3jINOJFFqavA9vzUjh8HyGZNzuj5OhBeZee03QmQLA2gfMBshDXxi6Y01VeA+QbrF
eSG3ngC8EQ7sVS2RYjran3ga8WGtBm3l8JJkyZSGUdeq6ed8b9MrUz6jMbQtOofyExjyEAUqyPy8
Bd5serx5AHwHMYcnizk9eTS9hDJJ8/ERYgIbgBg5nOyUGxa1O6Kww9Z1L9cZtJMV1565D6bwNF6g
j8Ropq1M+uvvY9rq9/XvAHQ3ap5Yyal99a7xuUTxHkOpq6e2v0ONDqqMe4cDGJortBxCqGggErW7
kptJGojtNMGSLSECMYKcM7uSyhR2ii7OoihXc3PQ2zmHCNDLUsoQqxPh7DgP0CfoGJPG3vTF7Apo
tGwbjTo2cGRL77BZelfl8WiTky2Syhy4TWrML3r/G5TFQjYjrrrLR3IWa6iBx9Ri3WuFGlAh2B3l
xk8zNhGNq07jS/7ljtYmPofp4BEmx9kM53YgfBCvneDMwI7g9HlLZ1dxeozIxE3+2skwGXMxHFv1
Wzto/42XpY35qcbsF/+lHPSnQEemvTeIbY3P3DOReAMhZ1xNEimi+NzgFZ3Q/WX/XDREkAan4bGs
xmca7OK0PoGWC4xVHq8FwgUJhQ3OjBO5H4c75CmmCrdhOyFC5fRQZ0xZwWEFNaVVeO9RmhWlxho5
mvmAaw1cm5jFKAvHAOROxBK2V+CiyXXvr0olu9A6Ya6tx2izeL1WIVJPTs9m4wFO8HNjsYsHPL4o
KOLmUJ9V2t5kG1NzO/1eWa4iA7IpElIybuA43FCegXsGcI9RUgJZ8vacxR/8+6bAWgCxZQS7RTMv
pFQoT+7KPQlFr6g/VADSxvKgefur+Po88dJp2Nh/VWGmsfz6AIDaqDZ0ip/OYd+Wh3r/o/eBpDLK
uw1xsua/X0hRlf+C2S7LrRo/twhQGFWlXLwwXMMmQQMaqnwfQhun5wxTWODUFJYI8v2+Qt3HTYdY
chKaF85shiGEnM/NyvhySY4OszxusYHwJEHk7PEtstTvEGaK+7GXm2zoUtokCUIEtMVSyr9YEQSM
RK3X5GtNy/zymYuQmwbpuRNygBYG79bVYv8VCrQsmxHx9YiFBnVLxJR179rJh2lsVC5Qk1hhxY8R
Bm0A0J37oIpqkICOv++zEytDyOtmwuZrFo1SW/g+YdqvckktHvkpm6d+nvGc8hbzQ8rcuu6TH5tw
v3YHy3K8CUe1fArp/+G5r3to1VsZIB9WmOnwALjAIo1C319//x24NCcNrKp/NMBreWOqIiooHCIC
+tFZtGLAKiv6wSEjZTn/oZ9WnggTiOEkV8vv4LUwOR16t+plk1x+/eshUepgKVh9RCZ5BrtVtApj
jTURjtfR13f+xkY5p8XexUyeRK6eEnjA+GmPOip+RWqpNFs4UHqo/upIpud0rGRtz4MrrdxGnYys
Heo9ed7oCTtbUPawutckP4VxEEpsTd/mDINjcl5R+uioId9BHZ/WhmP2X4uwSD4j/P7o6LVL2sm1
ioylIEUyuinukhIM8Kwec7gTYxhz9/iKteXz6H+HqzqXzOF0WZgiuSS4QTZhXV+ZfQ3fKSDb4wR4
ErphluGrHoYQfvOxvzo5ALJQp40aU4n5guPSz+3tnjZfC+CP7kqQ5rwowZw/KWNNOlOYzCeviyr7
CmNLCRCX7BJ21cAWb6xSMCeZZGF6SQl4KXpHOXDS/KqOyeRWez6EaSvRb62yOemLTQX5n1A5e68T
/u06wP+IB3B0SIlmcFs5Np3NSDG+lsFYafMEP/D5Uel45pmZJ1IHPDJIfHEMDS/n7arPw10XPaIY
cbDiSy/FgaeCNYg5SzkQVFtyJbRx2F5LybCLweDv8A6kL62h6olHqkSSrWN9ao+0niSb39KVHjjX
wz8ccd2L5U4RvtEF0Ris7S709ebfrdx/kXEggbfRHHd/n/SSMzOZyi3sy4d5PIY+OGAYqOZHMIJI
b2SddvfZALyqp0uk2f2uZTXbs3gSA8ltQ6miNX2Q8NnFjDdIx55bKwHgKgwo5uGncTfkheNgf1Mo
DC74gpcUM2J1iZgXvHB9JZV+nJA4GRkoWCIY5T5uY7j4UMVqob2Cb8PeUKDVSkJuqd+TQYLBm4+Y
ie+/SV7zefYN9PVTRMiis7FpXEOnREILWn98uMDEGLaJf3sIW+GBLCzOVM68QjW3hPxd8l5eft1g
NikozGUJi55AOfaSQtSLU6aXqS3oubV5EW1s2bjYWcw93IYFIB79DsJxxf6lle6SXx2uZCQJtXo5
S96PanttFPUISm2x/pA+0BeWjDSRavx7SqF3HeASbkEqEbao/ppo7YWbnyKxW9mLYMKcJML5nrSI
85PgthRSUPeJKUksCyMcY8zvP59dx1asskDYPcdyHbtuTcDNN0UYPNzEYcZ2Zoy1JTRMGl0O3JDA
HUBpezhXvGgAr3ZpKbyo2aW2vQwC2ehKaK3veBMLSg2KROhaXKH5mSGU4nY9maSGfYW80lFztK2q
VvBBD7myv9m448KARgjwvaiZzUpAhkQSIzIGfimvt9KIg+96J5XwTs788eX/S67F2tdezNuTmV54
MjiaU2nqr7xmlsUIxA3eabg++JYPNdm9dYogM2fM/a8jme8zeo+ioYm9dpardya2FFeuf6/HY6Kk
YB/qm5Q2k/Uxz+Dpj0Eo7YF3tFSnAkuj3gdg3kRJ06AehHFWJTca/q90RMOy7dlZ50HbBNMkJqnw
wdYobC52gkz85X1ADKo4/kw97ImWGII1e/XYeseaeFvygO4uVl7l1rHZ81DR2wkuDBzU4B9T4fm5
tKp5BaDCDP0ZRvpb4FYnE9YArWJi8gYRle9WY71O7XS84Vf8ksQLb6PyK8QiE7ETKtw0gdNeJKFy
Feol7O0QkYZ5+6nxOdNOEsRQa9eurzl1uItt4oZlNQzb2n1EUVlOf/dTzd3gQOcJteZj4K/709Pp
me2Gh2UjTxqZ1BCyYDtOfdFZ7118FfHkC59X/wzhHZAsBIrglgJGaVuRsJJ+WXis3uGank4sp+p3
NlUkROZu5PLsklAQt8xXdjL9KEWaKd6txzU30OUXmjpbeD4x5AawNCxdswtsX3cyBcd6PRp3JOGi
DM1H/b2c4qHBFTnGA0UkwBnhZkUoyNHNRsym9NNBwHnDdU5WxWOmmJiY0Y9UqBbO6n/yfxvJpM8u
VRWskbXSWm59wfdTJyPvZfTLfuLkU+l7NH2+PmPvwU9SptHHGEV9FO/hJucoSWDAfl2wUlynyFbZ
USwHKrGlectcn5dob3xyyLIdUWIaPkHaMuK+YTxszheXb1ECMtAm58CfjMtrGcvbbJflGHyHhrMU
Y5dR/ekJFw4xc8LCX36W+UMdqqai90UpbYwp92SfOGxSOccxdH4COB2q/T6KaceleK7iz1FlIhkP
adli2Q3ZsmAeHsHgcMcJ4W3sZ6joh9MTAqC3wNg2Hj11cziL2sDkfMv9t3rrC+8R0jcK4PPXclTW
FNLTSoZVjG81V3CtTQ4ex1iOQnyWpL7gRWI923W9Sbbj9uekYjJL2EEMnlAMV1k27suxFWrJIn1m
Jqu/sEhs4DDtmiZ2z87wNCq9BQj9clGvWAir4HiXBEQUMkcv1ORZtkRtQfuiMxW/NFd7pEAOYot3
FMLsfGeLTC1kSML+SGIrMlSWLyEeQIZA3jKXfMK3ocA0AYEzkrxMU6X+CU14DbyyTpotNsQIYQvm
PELzq0UyD0BYLfbnu4UlPuG6saBr9NkXKwA/sP23ElQtp5b1d7y/7uh+b62aIN8lkqoGaxeVPzl+
msNWc5NIBwHwk4TNUoYs6NkwoOYV6xHsaMOhhFRq+rRm3Z0A3Y5FkzgbAYdhAbRW/i0d9bruPhIh
KWMYpYzJ2gdRv80xRgVnMy38AY9eJQHrztzkN8mdnsaVry2xuep3Dia5Q5Ys0/eYEJStZMLRCijU
wJ3fccsHItebAY/zgY+pfLREI3fp5Npt2HFETWvb1im/ef8p2029TBA3ItpfbQtWPycjAnofuZA4
qMFn5WyLf3dmrCHH5AaiSlBzej2gKwaJ5ywfWscWfqtgmxyR/CxNINAJRR+d/Q/hMHCvLQJvIuQm
GjWT9mwdwtP7j+z34sgLZkTca1LtSh1WZkIs1xwT5WRxqigqhlYS3rNcNQevvtQ1e2OnPX3toFXt
0xXjvPmB3yFXFFPxDED9bGXXXe4lVA/AnlU/rxexqM804Xl4pBAuIsZ9/dZH9TkTg2dIjnAJ02Jd
Bs9GnDpChT6DQ/98Lc7TFazTfVDd3zWGxtM=
`protect end_protected
